`default_nettype none

module graphics
    #(
        parameter VGA_WIDTH = 640,
        parameter VGA_HEIGHT = 480,

        parameter H_FRONT_PORCH = 16,
        parameter H_SYNC_PULSE = 96,
        parameter H_BACK_PORCH = 48,

        parameter V_FRONT_PORCH = 10,
        parameter V_SYNC_PULSE = 2,
        parameter V_BACK_PORCH = 33
    )
    (
        input wire clk,
        input wire rst_n,

        output wire [7:0] vga_pmod
    );

    localparam X_PIXEL_BITS = $clog2(VGA_WIDTH);
    localparam Y_PIXEL_BITS = $clog2(VGA_HEIGHT);

    reg hsync;
    reg vsync;
    reg [1:0] red;
    reg [1:0] green;
    reg [1:0] blue;

    reg [X_PIXEL_BITS - 1 : 0] pixel_x;
    reg [Y_PIXEL_BITS - 1 : 0] pixel_y;

    assign vga_pmod = {hsync, blue[1], green[1], red[1], vsync, blue[0], green[0], red[0]};

    reg [203 : 0] bitmap [20 : 0];
    initial begin
        bitmap[0] = 204'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[1] = 204'b110100110100110100110100110100110100000000000000000000110100110100110100000000000000000000110100110100110100110100110100110100110100000000000000000000110100110100000000000000000000110100110100110100110100;
        bitmap[2] = 204'b110100110100110100110100110100110100000000010101010101000000110100000000010101010101000000110100110100110100110100110100110100000000010101010101000000110100000000010101010101000000110100110100110100110100;
        bitmap[3] = 204'b110100110100110100110100110100110100000000010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100;
        bitmap[4] = 204'b110100110100110100110100110100110100110100000000000000011011011011011011011011011011011011011011011011011011011011011011000000010101010101010101010101010101010101010101010101010101010101000000110100110100;
        bitmap[5] = 204'b110100110100110100110100110100110100110100000000011011011011011011110111110111110111110111110111110111110111110111000000010101010101010101000000000000000000000000000000000000000000010101010101000000110100;
        bitmap[6] = 204'b110100110100110100110100110100110100110100000000011011011011110111010011110111110111110111110111110111110111000000010101010111010111010101000000010101010101000000010101010101000000010101010111010111000000;
        bitmap[7] = 204'b110100110100110100110100110100000000000000000000011011110111110111110111110111110111010011110111110111110111000000010101010111010111010101010101010101010101010101010101010101010101010101010111010111000000;
        bitmap[8] = 204'b110100110100110100000000000000010101010101000000011011110111110111110111110111110111110111110111110111110111000000010101010101010101000000000000010101010101010101000000010101000000000000010101010101000000;
        bitmap[9] = 204'b110100110100000000010101010101010101010101000000011011110111010011110111110111110111110111110111110111110111000000010101010101010101111111000000010101010101010101010101010101111111000000010101010101000000;
        bitmap[10] = 204'b110100000000010101010101000000000000000000000000011011110111110111110111110111110111110111110111010011110111000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000;
        bitmap[11] = 204'b110100000000010101010101000000110100110100000000011011110111110111110111010011110111110111110111110111110111110111000000010101010101010101010101010101010101010101010101010101010101010101010101000000110100;
        bitmap[12] = 204'b110100110100000000000000110100110100110100000000011011110111110111110111110111110111110111110111110111110111110111000000010101010101010101010101000000000000000000000000010101010101010101010101000000110100;
        bitmap[13] = 204'b110100110100110100110100110100110100110100000000011011110111110111110111110111110111110111010011110111110111110111000000010101010101010101000000110111110111011011000000000000010101010101010101000000110100;
        bitmap[14] = 204'b110100110100110100110100110100110100110100000000011011110111110111110111110111110111110111110111110111110111110111000000010101010101000000110111110111110111011011000000110100000000010101010101000000110100;
        bitmap[15] = 204'b110100110100110100110100110100110100110100000000011011110111110111110111110111110111110111110111110111110111110111110111000000000000110111010011110111110111011011000000110100110100000000000000110100110100;
        bitmap[16] = 204'b110100110100110100110100110100110100110100000000011011110111110111010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011000000110100110100110100110100110100110100;
        bitmap[17] = 204'b110100110100110100110100110100110100110100000000011011011011110111110111110111110111110111110111010011110111110111010011110111110111110111110111110111011011011011000000110100110100110100110100110100110100;
        bitmap[18] = 204'b110100110100110100110100110100110100110100000000011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011000000110100110100110100110100110100110100;
        bitmap[19] = 204'b110100110100110100110100110100110100110100110100000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000110100110100110100110100110100110100110100;
        bitmap[20] = 204'b110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
    end         

    always @ (posedge clk) begin
        if (!rst_n) begin
            pixel_x <= {X_PIXEL_BITS{1'b0}};
            pixel_y <= {Y_PIXEL_BITS{1'b0}};
            hsync <= 1'b1;
            vsync <= 1'b1;
            red <= 2'd0;
            green <= 2'd0;
            blue <= 2'd0;
        end else begin
            if (pixel_x == VGA_WIDTH + H_FRONT_PORCH) begin
                hsync <= 1'b1;
            end
            if (pixel_x == VGA_WIDTH + H_FRONT_PORCH + H_SYNC_PULSE) begin
                hsync <= 1'b0;
            end

            if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH) begin
                vsync <= 1'b1;
            end
            if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH + V_SYNC_PULSE) begin
                vsync <= 1'b0;
            end

            if (pixel_x == VGA_WIDTH + H_BACK_PORCH + H_SYNC_PULSE + H_BACK_PORCH - 1) begin
                pixel_x <= {X_PIXEL_BITS{1'b0}};
                if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH + V_SYNC_PULSE + V_BACK_PORCH - 1) begin
                    pixel_y <= {Y_PIXEL_BITS{1'b0}};
                end else begin
                    pixel_y <= pixel_y + 1;
                end
            end else begin
                pixel_x <= pixel_x + 1;
            end

            if (pixel_x >= 100 && pixel_x < 100 + 34 * 8 && pixel_y > 100 && pixel_y < 100 + 21 * 8) begin
                {blue, green, red} <= bitmap[20 - (pixel_y - 100) / 8][(33 - (pixel_x - 100) / 8) * 6 + 5 -: 6];
            end else begin
                {red, green, blue} <= 6'b000111;
            end
            /*            
            if (pixel_x < VGA_WIDTH && pixel_y < VGA_HEIGHT) begin
                red <= random_value[1:0];
                green <= random_value[3:2];
                blue <= random_value[5:4];
            end else begin
                red <= 2'd0;
                green <= 2'd0;
                blue <= 2'd0;
            end
            */
        end
    end
endmodule

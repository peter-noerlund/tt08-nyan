// tt_um_vga_example

`default_nettype none

module tt_um_minesweeper
    (
        input wire [7:0] ui_in,
        output wire [7:0] uo_out,
        input wire [7:0] uio_in,
        output wire [7:0] uio_out,
        output wire [7:0] uio_oe,
        input wire ena,
        input wire clk,
        input wire rst_n
    );

    localparam HORI_WIDTH = 640;
    localparam HORI_FRONT_PORCH = 16;
    localparam HORI_SYNC_PULSE = 96;
    localparam HORI_BACK_PORCH = 48;

    localparam VERT_HEIGHT = 480;
    localparam VERT_FRONT_PORCH = 10;
    localparam VERT_SYNC_PULSE = 2;
    localparam VERT_BACK_PORCH = 33;
    
    localparam TILE_WIDTH = 32;
    localparam TILE_HEIGHT = 32;

    localparam HORI_TILES = HORI_WIDTH / TILE_WIDTH;
    localparam VERT_TILES = VERT_HEIGHT / TILE_HEIGHT;
    localparam TILE_COUNT = HORI_TILES * VERT_TILES;

    wire up;
    wire down;
    wire left;
    wire right;
    wire press;

    reg hsync;
    reg vsync;
    reg [1:0] red;
    reg [1:0] green;
    reg [1:0] blue;
    reg [9:0] x;
    reg [9:0] y;
    reg [4:0] cur_x;
    reg [4:0] cur_y;
    reg last_left;
    reg last_right;
    reg last_up;
    reg last_down;
    reg last_press;

    reg [TILE_COUNT - 1 : 0] state;
    reg [63:0] tile[31:0];
    reg [63:0] bomb[31:0];

    assign uio_oe = 8'b00000000;
    assign uio_out = 8'b00000000;
    assign uo_out = {hsync, blue[0], green[0], red[0], vsync, blue[1], green[1], red[1]};

    assign left = ui_in[0];
    assign right = ui_in[1];
    assign up = ui_in[2];
    assign down = ui_in[3];
    assign press = ui_in[4];

    always @ (posedge clk) begin
        if (!rst_n) begin
            x <= 10'd0;
            y <= 10'd0;
            hsync <= 1'b0;
            vsync <= 1'b0;
            red <= 2'd0;
            green <= 2'd0;
            blue <= 2'd0;
            cur_x <= 5'd0;
            cur_y <= 5'd0;
            last_left <= 1'b0;
            last_right <= 1'b0;
            last_up <= 1'b0;
            last_down <= 1'b0;
            last_press <= 1'b0;
            state <= {TILE_COUNT{1'b0}};
        end else begin
            if (x == HORI_WIDTH + HORI_FRONT_PORCH) begin
                hsync <= 1'b1;
            end
            if (x == HORI_WIDTH + HORI_FRONT_PORCH + HORI_SYNC_PULSE) begin
                hsync <= 1'b0;
            end
            if (y == VERT_HEIGHT + VERT_FRONT_PORCH) begin
                vsync <= 1'b1;
            end
            if (y == VERT_HEIGHT + VERT_FRONT_PORCH + VERT_SYNC_PULSE) begin
                vsync <= 1'b0;
            end

            if (x < HORI_WIDTH && y <= VERT_HEIGHT) begin
                if (x[9:5] == cur_x && y[9:5] == cur_y && (x[4:0] < 5'd2 || x[4:0] > 5'd29 || y[4:0] < 5'd2 || y[4:0] > 5'd29)) begin
                    red <= 2'd3;
                    green <= 2'd0;
                    blue <= 2'd0;
                end else if (state[y[9:5] * HORI_TILES + {5'd0, x[9:5]}] == 1'b0) begin
                    red <= tile[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                    green <= tile[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                    blue <= tile[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                end else begin
                    red <= bomb[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                    green <= bomb[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                    blue <= bomb[y & 31][(31 - x & 31) * 2 + 1 -: 2];
                end
            end else begin
                red <= 2'd0;
                green <= 2'd0;
                blue <= 2'd0;
            end

            if (x == HORI_WIDTH + HORI_FRONT_PORCH + HORI_SYNC_PULSE + HORI_BACK_PORCH - 1) begin
                x <= 10'd0;
                if (y == VERT_HEIGHT + VERT_FRONT_PORCH + VERT_SYNC_PULSE + VERT_BACK_PORCH - 1) begin
                    y <= 10'd0;
                end else begin
                    y <= y + 10'd1;
                end
            end else begin
                x <= x + 10'd1;
            end

            if (last_down && !down) begin
                cur_y <= cur_y + 5'd1;
            end else if (last_up && !up) begin
                cur_y <= cur_y - 5'd1;
            end

            if (last_left && !left) begin
                cur_x <= cur_x - 5'd1;
            end else if (last_right && !right) begin
                cur_x <= cur_x + 5'd1;
            end

            if (last_press && !press) begin
                state[{5'd0, cur_y} * HORI_TILES + {5'd0, cur_x}] <= 1'b1;
            end

            last_left <= left;
            last_up <= up;
            last_right <= right;
            last_down <= down;
            last_press <= press;
        end
    end

    initial begin
        tile[0]  = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        tile[1]  = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        tile[2]  = 64'b1111111111111111111111111111111111111111111111111111111111110101;
        tile[3]  = 64'b1111111111111111111111111111111111111111111111111111111111010101;
        tile[4]  = 64'b1111111111111111111111111111111111111111111111111111111101010101;
        tile[5]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[6]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[7]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[8]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[9]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[10] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[11] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[12] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[13] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[14] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[15] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[16] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[17] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[18] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[19] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[20] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[21] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[22] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[23] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[24] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[25] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[26] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[27] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[28] = 64'b1111110101010101010101010101010101010101010101010101010101010101;
        tile[29] = 64'b1111010101010101010101010101010101010101010101010101010101010101;
        tile[30] = 64'b1101010101010101010101010101010101010101010101010101010101010101;
        tile[31] = 64'b0101010101010101010101010101010101010101010101010101010101010101;

        bomb[0]  = 64'b01_01_01_01_01_01_01_01_01_01_01_0_101_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01;
        bomb[1]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[2]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[3]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[4]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[5]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[6]  = 64'b01_10_10_10_10_10_00_00_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_00_00_10_10_10_10_10_01;
        bomb[7]  = 64'b01_10_10_10_10_10_00_00_00_10_10_10_10_01_01_00_00_01_01_10_10_10_10_00_00_00_10_10_10_10_10_01;
        bomb[8]  = 64'b01_10_10_10_10_10_10_00_00_00_10_01_00_00_00_00_00_00_00_00_01_10_00_00_00_10_10_10_10_10_10_01;
        bomb[9]  = 64'b01_10_10_10_10_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_10_01;
        bomb[10] = 64'b01_10_10_10_10_10_10_10_10_00_00_00_00_01_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_10_10_01;
        bomb[11] = 64'b01_10_10_10_10_10_10_01_00_00_00_00_01_11_01_00_00_00_00_00_00_00_00_01_10_10_10_10_10_10_10_01;
        bomb[12] = 64'b01_10_10_10_10_10_10_00_00_00_00_01_11_11_01_00_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_01;
        bomb[13] = 64'b01_10_10_10_10_10_01_00_00_00_01_11_11_01_00_00_00_00_00_00_00_00_00_00_00_01_10_10_10_10_10_01;
        bomb[14] = 64'b01_10_10_10_10_10_01_00_00_00_00_01_01_00_00_00_00_00_00_00_00_00_00_00_00_01_10_10_10_10_10_01;
        bomb[15] = 64'b01_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_01;
        bomb[16] = 64'b01_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_01;
        bomb[17] = 64'b01_10_10_10_10_10_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_10_10_10_10_10_01;
        bomb[18] = 64'b01_10_10_10_10_10_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_10_10_10_10_10_01;
        bomb[19] = 64'b01_10_10_10_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_01;
        bomb[20] = 64'b01_10_10_10_10_10_10_01_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_01_10_10_10_10_10_10_10_01;
        bomb[21] = 64'b01_10_10_10_10_10_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_10_10_01;
        bomb[22]  = 64'b01_10_10_10_10_10_10_10_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_10_10_10_10_10_10_10_01;
        bomb[23]  = 64'b01_10_10_10_10_10_10_00_00_00_10_01_00_00_00_00_00_00_00_00_01_10_00_00_00_10_10_10_10_10_10_01;
        bomb[24]  = 64'b01_10_10_10_10_10_00_00_00_10_10_10_10_01_01_00_00_01_01_10_10_10_10_00_00_00_10_10_10_10_10_01;
        bomb[25]  = 64'b01_10_10_10_10_10_00_00_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_00_00_10_10_10_10_10_01;
        bomb[26]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[27]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_00_00_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[28]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[29]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[30]  = 64'b01_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_10_01;
        bomb[31]  = 64'b01_01_01_01_01_01_01_01_01_01_01_0_101_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01_01;
    end
endmodule

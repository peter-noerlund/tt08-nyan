// tt_um_vga_example

`timescale 1ns/1ps
`default_nettype none

module tt_um_minesweeper
    (
        input wire [7:0] ui_in,
        output wire [7:0] uo_out,
        input wire [7:0] uio_in,
        output wire [7:0] uio_out,
        output wire [7:0] uio_oe,
        input wire ena,
        input wire clk,
        input wire rst_n
    );

    localparam HORI_WIDTH = 640;
    localparam HORI_FRONT_PORCH = 16;
    localparam HORI_SYNC_PULSE = 96;
    localparam HORI_BACK_PORCH = 48;

    localparam VERT_HEIGHT = 480;
    localparam VERT_FRONT_PORCH = 10;
    localparam VERT_SYNC_PULSE = 2;
    localparam VERT_BACK_PORCH = 33;

    reg hsync;
    reg vsync;
    reg [1:0] color;
    reg [9:0] x;
    reg [9:0] y;

    reg [63:0] tile[31:0];

    assign uio_oe = 8'b00000000;
    assign uio_out = 8'b00000000;
    assign uo_out = {hsync, color[0], color[0], color[0], vsync, color[1], color[1], color[1]};

    always @ (posedge clk) begin
        if (!rst_n) begin
            x <= 10'd0;
            y <= 10'd0;
            hsync <= 1'b0;
            vsync <= 1'b0;
            color <= 2'd0;
        end else begin
            if (x == HORI_WIDTH + HORI_FRONT_PORCH) begin
                hsync <= 1'b1;
            end
            if (x == HORI_WIDTH + HORI_FRONT_PORCH + HORI_SYNC_PULSE) begin
                hsync <= 1'b0;
            end
            if (y == VERT_HEIGHT + VERT_FRONT_PORCH) begin
                vsync <= 1'b1;
            end
            if (y == VERT_HEIGHT + VERT_FRONT_PORCH + VERT_SYNC_PULSE) begin
                vsync <= 1'b0;
            end

            if (x < HORI_WIDTH && y <= HORI_WIDTH) begin
                color <= tile[y & 31][(31 - x & 31) * 2 + 1 -: 2];
            end

            if (x == HORI_WIDTH + HORI_FRONT_PORCH + HORI_SYNC_PULSE + HORI_BACK_PORCH - 1) begin
                x <= 10'd0;
                if (y == VERT_HEIGHT + VERT_FRONT_PORCH + VERT_SYNC_PULSE + VERT_BACK_PORCH - 1) begin
                    y <= 10'd0;
                end else begin
                    y <= y + 10'd1;
                end
            end else begin
                x <= x + 10'd1;
            end
        end
    end

    initial begin
        tile[0]  = 64'b1111111111111111111111111111111111111111111111111111111111111111;
        tile[1]  = 64'b1111111111111111111111111111111111111111111111111111111111111101;
        tile[2]  = 64'b1111111111111111111111111111111111111111111111111111111111110101;
        tile[3]  = 64'b1111111111111111111111111111111111111111111111111111111111010101;
        tile[4]  = 64'b1111111111111111111111111111111111111111111111111111111101010101;
        tile[5]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[6]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[7]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[8]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[9]  = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[10] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[11] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[12] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[13] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[14] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[15] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[16] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[17] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[18] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[19] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[20] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[21] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[22] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[23] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[24] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[25] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[26] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[27] = 64'b1111111110101010101010101010101010101010101010101010101001010101;
        tile[28] = 64'b1111110101010101010101010101010101010101010101010101010101010101;
        tile[29] = 64'b1111010101010101010101010101010101010101010101010101010101010101;
        tile[30] = 64'b1101010101010101010101010101010101010101010101010101010101010101;
        tile[31] = 64'b0101010101010101010101010101010101010101010101010101010101010101;
    end
endmodule
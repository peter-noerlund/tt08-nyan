initial begin
    // Section 1

    melody[0] = {B, LONG_NOTE};
    melody[1] = {LOW_F_SHARP, SHORT_NOTE};
    melody[2] = {LOW_G_SHARP, SHORT_NOTE};

    melody[3] = {B, LONG_NOTE};
    melody[4] = {LOW_F_SHARP, SHORT_NOTE};
    melody[5] = {LOW_G_SHARP, SHORT_NOTE};

    melody[6] = {B, SHORT_NOTE};
    melody[7] = {C_SHARP, SHORT_NOTE};
    melody[8] = {D_SHARP, SHORT_NOTE};
    melody[9] = {B, SHORT_NOTE};

    melody[10] = {E, SHORT_NOTE};
    melody[11] = {D_SHARP, SHORT_NOTE};
    melody[12] = {E, SHORT_NOTE};
    melody[13] = {F_SHARP, SHORT_NOTE};

    // Section 2

    melody[14] = {B, LONG_NOTE};
    melody[15] = {B, LONG_NOTE};

    melody[16] = {LOW_F_SHARP, SHORT_NOTE};
    melody[17] = {LOW_G_SHARP, SHORT_NOTE};
    melody[18] = {B, SHORT_NOTE};
    melody[19] = {LOW_F_SHARP, SHORT_NOTE};

    melody[20] = {E, SHORT_NOTE};
    melody[21] = {D_SHARP, SHORT_NOTE};
    melody[22] = {C_SHARP, SHORT_NOTE};
    melody[23] = {B, SHORT_NOTE};

    melody[24] = {LOW_F_SHARP, SHORT_NOTE};
    melody[25] = {LOW_D_SHARP, SHORT_NOTE};
    melody[26] = {LOW_E, SHORT_NOTE};
    melody[27] = {LOW_F_SHARP, SHORT_NOTE};

    // Section 3

    melody[28] = {B, LONG_NOTE};
    melody[29] = {LOW_F_SHARP, SHORT_NOTE};
    melody[30] = {LOW_G_SHARP, SHORT_NOTE};

    melody[31] = {B, LONG_NOTE};
    melody[32] = {LOW_F_SHARP, SHORT_NOTE};
    melody[33] = {LOW_G_SHARP, SHORT_NOTE};

    melody[34] = {B, SHORT_NOTE};
    melody[35] = {B, SHORT_NOTE};
    melody[36] = {C_SHARP, SHORT_NOTE};
    melody[37] = {D_SHARP, SHORT_NOTE};

    melody[38] = {B, SHORT_NOTE};
    melody[39] = {LOW_F_SHARP, SHORT_NOTE};
    melody[40] = {LOW_G_SHARP, SHORT_NOTE};
    melody[41] = {LOW_F_SHARP, SHORT_NOTE};

    // Section 4
    
    melody[42] = {B, LONG_NOTE};
    melody[43] = {B, SHORT_NOTE};
    melody[44] = {LOW_A_SHARP, SHORT_NOTE};

    melody[45] = {B, SHORT_NOTE};
    melody[46] = {LOW_F_SHARP, SHORT_NOTE};
    melody[47] = {LOW_G_SHARP, SHORT_NOTE};
    melody[48] = {B, SHORT_NOTE};

    melody[49] = {E, SHORT_NOTE};
    melody[50] = {D_SHARP, SHORT_NOTE};
    melody[51] = {E, SHORT_NOTE};
    melody[52] = {F_SHARP, SHORT_NOTE};

    melody[53] = {B, LONG_NOTE};
    melody[54] = {LOW_A_SHARP, LONG_NOTE};

    // Section 5

    melody[55] = {B, LONG_NOTE};
    melody[56] = {LOW_F_SHARP, SHORT_NOTE};
    melody[57] = {LOW_G_SHARP, SHORT_NOTE};

    melody[58] = {B, LONG_NOTE};
    melody[59] = {LOW_F_SHARP, SHORT_NOTE};
    melody[60] = {LOW_G_SHARP, SHORT_NOTE};

    melody[61] = {B, SHORT_NOTE};
    melody[62] = {C_SHARP, SHORT_NOTE};
    melody[63] = {D_SHARP, SHORT_NOTE};
    melody[64] = {B, SHORT_NOTE};

    melody[65] = {E, SHORT_NOTE};
    melody[66] = {D_SHARP, SHORT_NOTE};
    melody[67] = {E, SHORT_NOTE};
    melody[68] = {F_SHARP, SHORT_NOTE};

    // Section 6

    melody[69] = {B, LONG_NOTE};
    melody[70] = {B, LONG_NOTE};

    melody[71] = {LOW_F_SHARP, SHORT_NOTE};
    melody[72] = {LOW_G_SHARP, SHORT_NOTE};
    melody[73] = {B, SHORT_NOTE};
    melody[74] = {LOW_F_SHARP, SHORT_NOTE};

    melody[75] = {E, SHORT_NOTE};
    melody[76] = {D_SHARP, SHORT_NOTE};
    melody[77] = {C_SHARP, SHORT_NOTE};
    melody[78] = {B, SHORT_NOTE};

    melody[79] = {LOW_F_SHARP, SHORT_NOTE};
    melody[80] = {LOW_D_SHARP, SHORT_NOTE};
    melody[81] = {LOW_E, SHORT_NOTE};
    melody[82] = {LOW_F_SHARP, SHORT_NOTE};

    // Section 7

    melody[83] = {B, LONG_NOTE};
    melody[84] = {LOW_F_SHARP, SHORT_NOTE};
    melody[85] = {LOW_G_SHARP, SHORT_NOTE};

    melody[86] = {B, LONG_NOTE};
    melody[87] = {LOW_F_SHARP, SHORT_NOTE};
    melody[88] = {LOW_G_SHARP, SHORT_NOTE};

    melody[89] = {B, SHORT_NOTE};
    melody[90] = {B, SHORT_NOTE};
    melody[91] = {C_SHARP, SHORT_NOTE};
    melody[92] = {D_SHARP, SHORT_NOTE};

    melody[93] = {B, SHORT_NOTE};
    melody[94] = {LOW_F_SHARP, SHORT_NOTE};
    melody[95] = {LOW_G_SHARP, SHORT_NOTE};
    melody[96] = {LOW_F_SHARP, SHORT_NOTE};

    // Section 8
    
    melody[97] = {B, LONG_NOTE};
    melody[98] = {B, SHORT_NOTE};
    melody[99] = {LOW_A_SHARP, SHORT_NOTE};

    melody[100] = {B, SHORT_NOTE};
    melody[101] = {LOW_F_SHARP, SHORT_NOTE};
    melody[102] = {LOW_G_SHARP, SHORT_NOTE};
    melody[103] = {B, SHORT_NOTE};

    melody[104] = {E, SHORT_NOTE};
    melody[105] = {D_SHARP, SHORT_NOTE};
    melody[106] = {E, SHORT_NOTE};
    melody[107] = {F_SHARP, SHORT_NOTE};

    melody[108] = {B, LONG_NOTE};
    melody[109] = {C_SHARP, LONG_NOTE};

    // Section 9

    melody[110] = {F_SHARP, LONG_NOTE};
    melody[111] = {G_SHARP, LONG_NOTE};
    
    melody[112] = {D, SHORT_NOTE};
    melody[113] = {D_SHARP, LONG_NOTE};
    melody[114] = {B, SHORT_NOTE};
    
    melody[115] = {D, SHORT_NOTE};
    melody[116] = {C_SHARP, SHORT_NOTE};
    melody[117] = {B, LONG_NOTE};
    
    melody[118] = {B, LONG_NOTE};
    melody[119] = {C_SHARP, LONG_NOTE};
    
    // Section 10

    melody[120] = {D, LONG_NOTE};
    melody[121] = {D, SHORT_NOTE};
    melody[122] = {C_SHARP, SHORT_NOTE};
    
    melody[123] = {B, SHORT_NOTE};
    melody[124] = {C_SHARP, SHORT_NOTE};
    melody[125] = {D_SHARP, SHORT_NOTE};
    melody[126] = {F_SHARP, SHORT_NOTE};
    
    melody[127] = {G_SHARP, SHORT_NOTE};
    melody[128] = {D_SHARP, SHORT_NOTE};
    melody[129] = {F_SHARP, SHORT_NOTE};
    melody[130] = {C_SHARP, SHORT_NOTE};
    
    melody[131] = {D, SHORT_NOTE};
    melody[132] = {B, SHORT_NOTE};
    melody[133] = {C_SHARP, SHORT_NOTE};
    melody[134] = {B, SHORT_NOTE};
    
    // Section 11
    
    melody[135] = {D_SHARP, LONG_NOTE};
    melody[136] = {F_SHARP, LONG_NOTE};
    
    melody[137] = {G_SHARP, SHORT_NOTE};
    melody[138] = {G_SHARP, SHORT_NOTE};
    melody[139] = {F_SHARP, SHORT_NOTE};
    melody[140] = {C_SHARP, SHORT_NOTE};
    
    melody[141] = {D_SHARP, SHORT_NOTE};
    melody[142] = {B, SHORT_NOTE};
    melody[143] = {D, SHORT_NOTE};
    melody[144] = {D_SHARP, SHORT_NOTE};
    
    melody[145] = {D, SHORT_NOTE};
    melody[146] = {C_SHARP, SHORT_NOTE};
    melody[147] = {B, SHORT_NOTE};
    melody[148] = {C_SHARP, SHORT_NOTE};
    
    // Section 12
    
    melody[149] = {D, LONG_NOTE};
    melody[150] = {B, SHORT_NOTE};
    melody[151] = {C_SHARP, SHORT_NOTE};
    
    melody[152] = {D_SHARP, SHORT_NOTE};
    melody[153] = {F_SHARP, SHORT_NOTE};
    melody[154] = {C_SHARP, SHORT_NOTE};
    melody[155] = {D, SHORT_NOTE};
    
    melody[156] = {C_SHARP, SHORT_NOTE};
    melody[157] = {B, SHORT_NOTE};
    melody[158] = {C_SHARP, LONG_NOTE};

    melody[159] = {B, LONG_NOTE};
    melody[160] = {C_SHARP, LONG_NOTE};
    
    // Section 13
    
    melody[161] = {F_SHARP, LONG_NOTE};
    melody[162] = {G_SHARP, LONG_NOTE};
    
    melody[163] = {D, SHORT_NOTE};
    melody[164] = {D_SHARP, LONG_NOTE};
    melody[165] = {B, SHORT_NOTE};
    
    melody[166] = {D, SHORT_NOTE};
    melody[167] = {C_SHARP, SHORT_NOTE};
    melody[168] = {B, LONG_NOTE};
    
    melody[169] = {B, LONG_NOTE};
    melody[170] = {C_SHARP, LONG_NOTE};
    
    // Section 14
    
    melody[171] = {D, LONG_NOTE};
    melody[172] = {D, SHORT_NOTE};
    melody[173] = {C_SHARP, SHORT_NOTE};
    
    melody[174] = {B, SHORT_NOTE};
    melody[175] = {C_SHARP, SHORT_NOTE};
    melody[176] = {D_SHARP, SHORT_NOTE};
    melody[177] = {F_SHARP, SHORT_NOTE};
    
    melody[178] = {G_SHARP, SHORT_NOTE};
    melody[179] = {D_SHARP, SHORT_NOTE};
    melody[180] = {F_SHARP, SHORT_NOTE};
    melody[181] = {C_SHARP, SHORT_NOTE};
    
    melody[182] = {D, SHORT_NOTE};
    melody[183] = {B, SHORT_NOTE};
    melody[184] = {C_SHARP, SHORT_NOTE};
    melody[185] = {B, SHORT_NOTE};
    
    // Section 15
    
    melody[186] = {D_SHARP, LONG_NOTE};
    melody[187] = {F_SHARP, LONG_NOTE};
    
    melody[188] = {G_SHARP, SHORT_NOTE};
    melody[189] = {G_SHARP, SHORT_NOTE};
    melody[190] = {F_SHARP, SHORT_NOTE};
    melody[191] = {C_SHARP, SHORT_NOTE};
    
    melody[192] = {D_SHARP, SHORT_NOTE};
    melody[193] = {B, SHORT_NOTE};
    melody[194] = {D, SHORT_NOTE};
    melody[195] = {D_SHARP, SHORT_NOTE};
    
    melody[196] = {D, SHORT_NOTE};
    melody[197] = {C_SHARP, SHORT_NOTE};
    melody[198] = {B, SHORT_NOTE};
    melody[199] = {C_SHARP, SHORT_NOTE};
    
    // Section 16
    
    melody[200] = {D, LONG_NOTE};
    melody[201] = {B, SHORT_NOTE};
    melody[202] = {C_SHARP, SHORT_NOTE};
    
    melody[203] = {D_SHARP, SHORT_NOTE};
    melody[204] = {F_SHARP, SHORT_NOTE};
    melody[205] = {C_SHARP, SHORT_NOTE};
    melody[206] = {D, SHORT_NOTE};
    
    melody[207] = {C_SHARP, SHORT_NOTE};
    melody[208] = {B, SHORT_NOTE};
    melody[209] = {C_SHARP, LONG_NOTE};
    
    melody[210] = {B, LONG_NOTE};
    melody[211] = {B, LONG_NOTE};
end

reg [4:0] frame0[31:0][47:0];
initial begin
    frame0[0][0] = 5'd0;
    frame0[1][0] = 5'd0;
    frame0[2][0] = 5'd0;
    frame0[3][0] = 5'd0;
    frame0[4][0] = 5'd0;
    frame0[5][0] = 5'd0;
    frame0[6][0] = 5'd0;
    frame0[7][0] = 5'd0;
    frame0[8][0] = 5'd0;
    frame0[9][0] = 5'd0;
    frame0[10][0] = 5'd0;
    frame0[11][0] = 5'd0;
    frame0[12][0] = 5'd0;
    frame0[13][0] = 5'd0;
    frame0[14][0] = 5'd0;
    frame0[15][0] = 5'd0;
    frame0[16][0] = 5'd0;
    frame0[17][0] = 5'd0;
    frame0[18][0] = 5'd0;
    frame0[19][0] = 5'd0;
    frame0[20][0] = 5'd0;
    frame0[21][0] = 5'd0;
    frame0[22][0] = 5'd0;
    frame0[23][0] = 5'd0;
    frame0[24][0] = 5'd0;
    frame0[25][0] = 5'd0;
    frame0[26][0] = 5'd0;
    frame0[27][0] = 5'd0;
    frame0[28][0] = 5'd0;
    frame0[29][0] = 5'd0;
    frame0[30][0] = 5'd0;
    frame0[31][0] = 5'd0;
    frame0[0][1] = 5'd0;
    frame0[1][1] = 5'd0;
    frame0[2][1] = 5'd0;
    frame0[3][1] = 5'd0;
    frame0[4][1] = 5'd0;
    frame0[5][1] = 5'd0;
    frame0[6][1] = 5'd0;
    frame0[7][1] = 5'd0;
    frame0[8][1] = 5'd0;
    frame0[9][1] = 5'd0;
    frame0[10][1] = 5'd0;
    frame0[11][1] = 5'd0;
    frame0[12][1] = 5'd0;
    frame0[13][1] = 5'd0;
    frame0[14][1] = 5'd0;
    frame0[15][1] = 5'd0;
    frame0[16][1] = 5'd0;
    frame0[17][1] = 5'd0;
    frame0[18][1] = 5'd0;
    frame0[19][1] = 5'd0;
    frame0[20][1] = 5'd0;
    frame0[21][1] = 5'd0;
    frame0[22][1] = 5'd0;
    frame0[23][1] = 5'd0;
    frame0[24][1] = 5'd0;
    frame0[25][1] = 5'd0;
    frame0[26][1] = 5'd0;
    frame0[27][1] = 5'd0;
    frame0[28][1] = 5'd0;
    frame0[29][1] = 5'd0;
    frame0[30][1] = 5'd0;
    frame0[31][1] = 5'd0;
    frame0[0][2] = 5'd0;
    frame0[1][2] = 5'd0;
    frame0[2][2] = 5'd0;
    frame0[3][2] = 5'd0;
    frame0[4][2] = 5'd0;
    frame0[5][2] = 5'd0;
    frame0[6][2] = 5'd0;
    frame0[7][2] = 5'd0;
    frame0[8][2] = 5'd0;
    frame0[9][2] = 5'd0;
    frame0[10][2] = 5'd0;
    frame0[11][2] = 5'd0;
    frame0[12][2] = 5'd0;
    frame0[13][2] = 5'd0;
    frame0[14][2] = 5'd0;
    frame0[15][2] = 5'd0;
    frame0[16][2] = 5'd0;
    frame0[17][2] = 5'd0;
    frame0[18][2] = 5'd0;
    frame0[19][2] = 5'd0;
    frame0[20][2] = 5'd0;
    frame0[21][2] = 5'd0;
    frame0[22][2] = 5'd0;
    frame0[23][2] = 5'd0;
    frame0[24][2] = 5'd0;
    frame0[25][2] = 5'd0;
    frame0[26][2] = 5'd0;
    frame0[27][2] = 5'd0;
    frame0[28][2] = 5'd0;
    frame0[29][2] = 5'd0;
    frame0[30][2] = 5'd0;
    frame0[31][2] = 5'd0;
    frame0[0][3] = 5'd0;
    frame0[1][3] = 5'd0;
    frame0[2][3] = 5'd0;
    frame0[3][3] = 5'd0;
    frame0[4][3] = 5'd0;
    frame0[5][3] = 5'd0;
    frame0[6][3] = 5'd0;
    frame0[7][3] = 5'd0;
    frame0[8][3] = 5'd0;
    frame0[9][3] = 5'd0;
    frame0[10][3] = 5'd0;
    frame0[11][3] = 5'd0;
    frame0[12][3] = 5'd0;
    frame0[13][3] = 5'd0;
    frame0[14][3] = 5'd0;
    frame0[15][3] = 5'd0;
    frame0[16][3] = 5'd0;
    frame0[17][3] = 5'd0;
    frame0[18][3] = 5'd0;
    frame0[19][3] = 5'd0;
    frame0[20][3] = 5'd0;
    frame0[21][3] = 5'd0;
    frame0[22][3] = 5'd0;
    frame0[23][3] = 5'd0;
    frame0[24][3] = 5'd0;
    frame0[25][3] = 5'd0;
    frame0[26][3] = 5'd0;
    frame0[27][3] = 5'd0;
    frame0[28][3] = 5'd0;
    frame0[29][3] = 5'd0;
    frame0[30][3] = 5'd0;
    frame0[31][3] = 5'd0;
    frame0[0][4] = 5'd0;
    frame0[1][4] = 5'd0;
    frame0[2][4] = 5'd0;
    frame0[3][4] = 5'd0;
    frame0[4][4] = 5'd0;
    frame0[5][4] = 5'd0;
    frame0[6][4] = 5'd0;
    frame0[7][4] = 5'd0;
    frame0[8][4] = 5'd0;
    frame0[9][4] = 5'd0;
    frame0[10][4] = 5'd0;
    frame0[11][4] = 5'd0;
    frame0[12][4] = 5'd0;
    frame0[13][4] = 5'd0;
    frame0[14][4] = 5'd0;
    frame0[15][4] = 5'd0;
    frame0[16][4] = 5'd0;
    frame0[17][4] = 5'd0;
    frame0[18][4] = 5'd0;
    frame0[19][4] = 5'd0;
    frame0[20][4] = 5'd0;
    frame0[21][4] = 5'd0;
    frame0[22][4] = 5'd0;
    frame0[23][4] = 5'd0;
    frame0[24][4] = 5'd0;
    frame0[25][4] = 5'd0;
    frame0[26][4] = 5'd0;
    frame0[27][4] = 5'd0;
    frame0[28][4] = 5'd0;
    frame0[29][4] = 5'd0;
    frame0[30][4] = 5'd0;
    frame0[31][4] = 5'd0;
    frame0[0][5] = 5'd0;
    frame0[1][5] = 5'd0;
    frame0[2][5] = 5'd0;
    frame0[3][5] = 5'd0;
    frame0[4][5] = 5'd0;
    frame0[5][5] = 5'd0;
    frame0[6][5] = 5'd0;
    frame0[7][5] = 5'd0;
    frame0[8][5] = 5'd0;
    frame0[9][5] = 5'd0;
    frame0[10][5] = 5'd0;
    frame0[11][5] = 5'd0;
    frame0[12][5] = 5'd0;
    frame0[13][5] = 5'd0;
    frame0[14][5] = 5'd0;
    frame0[15][5] = 5'd0;
    frame0[16][5] = 5'd0;
    frame0[17][5] = 5'd0;
    frame0[18][5] = 5'd0;
    frame0[19][5] = 5'd0;
    frame0[20][5] = 5'd0;
    frame0[21][5] = 5'd0;
    frame0[22][5] = 5'd0;
    frame0[23][5] = 5'd0;
    frame0[24][5] = 5'd0;
    frame0[25][5] = 5'd0;
    frame0[26][5] = 5'd0;
    frame0[27][5] = 5'd0;
    frame0[28][5] = 5'd0;
    frame0[29][5] = 5'd0;
    frame0[30][5] = 5'd0;
    frame0[31][5] = 5'd0;
    frame0[0][6] = 5'd0;
    frame0[1][6] = 5'd0;
    frame0[2][6] = 5'd0;
    frame0[3][6] = 5'd0;
    frame0[4][6] = 5'd0;
    frame0[5][6] = 5'd0;
    frame0[6][6] = 5'd0;
    frame0[7][6] = 5'd0;
    frame0[8][6] = 5'd0;
    frame0[9][6] = 5'd0;
    frame0[10][6] = 5'd0;
    frame0[11][6] = 5'd0;
    frame0[12][6] = 5'd0;
    frame0[13][6] = 5'd0;
    frame0[14][6] = 5'd0;
    frame0[15][6] = 5'd0;
    frame0[16][6] = 5'd0;
    frame0[17][6] = 5'd0;
    frame0[18][6] = 5'd0;
    frame0[19][6] = 5'd0;
    frame0[20][6] = 5'd0;
    frame0[21][6] = 5'd0;
    frame0[22][6] = 5'd0;
    frame0[23][6] = 5'd0;
    frame0[24][6] = 5'd0;
    frame0[25][6] = 5'd0;
    frame0[26][6] = 5'd0;
    frame0[27][6] = 5'd0;
    frame0[28][6] = 5'd0;
    frame0[29][6] = 5'd0;
    frame0[30][6] = 5'd0;
    frame0[31][6] = 5'd0;
    frame0[0][7] = 5'd0;
    frame0[1][7] = 5'd0;
    frame0[2][7] = 5'd0;
    frame0[3][7] = 5'd0;
    frame0[4][7] = 5'd0;
    frame0[5][7] = 5'd0;
    frame0[6][7] = 5'd0;
    frame0[7][7] = 5'd0;
    frame0[8][7] = 5'd0;
    frame0[9][7] = 5'd0;
    frame0[10][7] = 5'd0;
    frame0[11][7] = 5'd0;
    frame0[12][7] = 5'd0;
    frame0[13][7] = 5'd0;
    frame0[14][7] = 5'd0;
    frame0[15][7] = 5'd0;
    frame0[16][7] = 5'd0;
    frame0[17][7] = 5'd0;
    frame0[18][7] = 5'd0;
    frame0[19][7] = 5'd0;
    frame0[20][7] = 5'd0;
    frame0[21][7] = 5'd0;
    frame0[22][7] = 5'd0;
    frame0[23][7] = 5'd0;
    frame0[24][7] = 5'd0;
    frame0[25][7] = 5'd0;
    frame0[26][7] = 5'd0;
    frame0[27][7] = 5'd0;
    frame0[28][7] = 5'd0;
    frame0[29][7] = 5'd0;
    frame0[30][7] = 5'd0;
    frame0[31][7] = 5'd0;
    frame0[0][8] = 5'd0;
    frame0[1][8] = 5'd0;
    frame0[2][8] = 5'd0;
    frame0[3][8] = 5'd0;
    frame0[4][8] = 5'd0;
    frame0[5][8] = 5'd0;
    frame0[6][8] = 5'd0;
    frame0[7][8] = 5'd0;
    frame0[8][8] = 5'd0;
    frame0[9][8] = 5'd0;
    frame0[10][8] = 5'd0;
    frame0[11][8] = 5'd0;
    frame0[12][8] = 5'd0;
    frame0[13][8] = 5'd0;
    frame0[14][8] = 5'd0;
    frame0[15][8] = 5'd0;
    frame0[16][8] = 5'd0;
    frame0[17][8] = 5'd0;
    frame0[18][8] = 5'd0;
    frame0[19][8] = 5'd0;
    frame0[20][8] = 5'd0;
    frame0[21][8] = 5'd0;
    frame0[22][8] = 5'd0;
    frame0[23][8] = 5'd0;
    frame0[24][8] = 5'd0;
    frame0[25][8] = 5'd0;
    frame0[26][8] = 5'd0;
    frame0[27][8] = 5'd0;
    frame0[28][8] = 5'd0;
    frame0[29][8] = 5'd0;
    frame0[30][8] = 5'd0;
    frame0[31][8] = 5'd0;
    frame0[0][9] = 5'd0;
    frame0[1][9] = 5'd0;
    frame0[2][9] = 5'd0;
    frame0[3][9] = 5'd0;
    frame0[4][9] = 5'd0;
    frame0[5][9] = 5'd0;
    frame0[6][9] = 5'd0;
    frame0[7][9] = 5'd0;
    frame0[8][9] = 5'd0;
    frame0[9][9] = 5'd0;
    frame0[10][9] = 5'd0;
    frame0[11][9] = 5'd0;
    frame0[12][9] = 5'd0;
    frame0[13][9] = 5'd0;
    frame0[14][9] = 5'd0;
    frame0[15][9] = 5'd0;
    frame0[16][9] = 5'd0;
    frame0[17][9] = 5'd0;
    frame0[18][9] = 5'd0;
    frame0[19][9] = 5'd0;
    frame0[20][9] = 5'd0;
    frame0[21][9] = 5'd0;
    frame0[22][9] = 5'd0;
    frame0[23][9] = 5'd0;
    frame0[24][9] = 5'd0;
    frame0[25][9] = 5'd0;
    frame0[26][9] = 5'd0;
    frame0[27][9] = 5'd0;
    frame0[28][9] = 5'd0;
    frame0[29][9] = 5'd0;
    frame0[30][9] = 5'd0;
    frame0[31][9] = 5'd0;
    frame0[0][10] = 5'd0;
    frame0[1][10] = 5'd0;
    frame0[2][10] = 5'd0;
    frame0[3][10] = 5'd0;
    frame0[4][10] = 5'd0;
    frame0[5][10] = 5'd0;
    frame0[6][10] = 5'd0;
    frame0[7][10] = 5'd0;
    frame0[8][10] = 5'd0;
    frame0[9][10] = 5'd0;
    frame0[10][10] = 5'd0;
    frame0[11][10] = 5'd0;
    frame0[12][10] = 5'd0;
    frame0[13][10] = 5'd0;
    frame0[14][10] = 5'd0;
    frame0[15][10] = 5'd0;
    frame0[16][10] = 5'd0;
    frame0[17][10] = 5'd0;
    frame0[18][10] = 5'd0;
    frame0[19][10] = 5'd0;
    frame0[20][10] = 5'd0;
    frame0[21][10] = 5'd0;
    frame0[22][10] = 5'd0;
    frame0[23][10] = 5'd0;
    frame0[24][10] = 5'd0;
    frame0[25][10] = 5'd0;
    frame0[26][10] = 5'd0;
    frame0[27][10] = 5'd0;
    frame0[28][10] = 5'd0;
    frame0[29][10] = 5'd0;
    frame0[30][10] = 5'd0;
    frame0[31][10] = 5'd0;
    frame0[0][11] = 5'd0;
    frame0[1][11] = 5'd0;
    frame0[2][11] = 5'd0;
    frame0[3][11] = 5'd0;
    frame0[4][11] = 5'd0;
    frame0[5][11] = 5'd0;
    frame0[6][11] = 5'd0;
    frame0[7][11] = 5'd0;
    frame0[8][11] = 5'd0;
    frame0[9][11] = 5'd0;
    frame0[10][11] = 5'd0;
    frame0[11][11] = 5'd0;
    frame0[12][11] = 5'd0;
    frame0[13][11] = 5'd0;
    frame0[14][11] = 5'd0;
    frame0[15][11] = 5'd0;
    frame0[16][11] = 5'd0;
    frame0[17][11] = 5'd0;
    frame0[18][11] = 5'd0;
    frame0[19][11] = 5'd0;
    frame0[20][11] = 5'd0;
    frame0[21][11] = 5'd0;
    frame0[22][11] = 5'd0;
    frame0[23][11] = 5'd0;
    frame0[24][11] = 5'd0;
    frame0[25][11] = 5'd0;
    frame0[26][11] = 5'd0;
    frame0[27][11] = 5'd0;
    frame0[28][11] = 5'd0;
    frame0[29][11] = 5'd0;
    frame0[30][11] = 5'd0;
    frame0[31][11] = 5'd0;
    frame0[0][12] = 5'd0;
    frame0[1][12] = 5'd0;
    frame0[2][12] = 5'd0;
    frame0[3][12] = 5'd0;
    frame0[4][12] = 5'd0;
    frame0[5][12] = 5'd0;
    frame0[6][12] = 5'd0;
    frame0[7][12] = 5'd0;
    frame0[8][12] = 5'd0;
    frame0[9][12] = 5'd0;
    frame0[10][12] = 5'd0;
    frame0[11][12] = 5'd0;
    frame0[12][12] = 5'd0;
    frame0[13][12] = 5'd0;
    frame0[14][12] = 5'd0;
    frame0[15][12] = 5'd0;
    frame0[16][12] = 5'd0;
    frame0[17][12] = 5'd0;
    frame0[18][12] = 5'd0;
    frame0[19][12] = 5'd0;
    frame0[20][12] = 5'd0;
    frame0[21][12] = 5'd0;
    frame0[22][12] = 5'd0;
    frame0[23][12] = 5'd0;
    frame0[24][12] = 5'd0;
    frame0[25][12] = 5'd0;
    frame0[26][12] = 5'd0;
    frame0[27][12] = 5'd0;
    frame0[28][12] = 5'd0;
    frame0[29][12] = 5'd0;
    frame0[30][12] = 5'd0;
    frame0[31][12] = 5'd0;
    frame0[0][13] = 5'd0;
    frame0[1][13] = 5'd0;
    frame0[2][13] = 5'd0;
    frame0[3][13] = 5'd0;
    frame0[4][13] = 5'd0;
    frame0[5][13] = 5'd0;
    frame0[6][13] = 5'd0;
    frame0[7][13] = 5'd0;
    frame0[8][13] = 5'd0;
    frame0[9][13] = 5'd0;
    frame0[10][13] = 5'd0;
    frame0[11][13] = 5'd0;
    frame0[12][13] = 5'd0;
    frame0[13][13] = 5'd0;
    frame0[14][13] = 5'd0;
    frame0[15][13] = 5'd0;
    frame0[16][13] = 5'd0;
    frame0[17][13] = 5'd0;
    frame0[18][13] = 5'd0;
    frame0[19][13] = 5'd0;
    frame0[20][13] = 5'd0;
    frame0[21][13] = 5'd0;
    frame0[22][13] = 5'd0;
    frame0[23][13] = 5'd0;
    frame0[24][13] = 5'd0;
    frame0[25][13] = 5'd0;
    frame0[26][13] = 5'd0;
    frame0[27][13] = 5'd0;
    frame0[28][13] = 5'd0;
    frame0[29][13] = 5'd0;
    frame0[30][13] = 5'd0;
    frame0[31][13] = 5'd0;
    frame0[0][14] = 5'd0;
    frame0[1][14] = 5'd0;
    frame0[2][14] = 5'd0;
    frame0[3][14] = 5'd0;
    frame0[4][14] = 5'd0;
    frame0[5][14] = 5'd0;
    frame0[6][14] = 5'd0;
    frame0[7][14] = 5'd0;
    frame0[8][14] = 5'd0;
    frame0[9][14] = 5'd0;
    frame0[10][14] = 5'd0;
    frame0[11][14] = 5'd0;
    frame0[12][14] = 5'd0;
    frame0[13][14] = 5'd0;
    frame0[14][14] = 5'd0;
    frame0[15][14] = 5'd0;
    frame0[16][14] = 5'd0;
    frame0[17][14] = 5'd0;
    frame0[18][14] = 5'd0;
    frame0[19][14] = 5'd0;
    frame0[20][14] = 5'd0;
    frame0[21][14] = 5'd0;
    frame0[22][14] = 5'd0;
    frame0[23][14] = 5'd0;
    frame0[24][14] = 5'd0;
    frame0[25][14] = 5'd0;
    frame0[26][14] = 5'd0;
    frame0[27][14] = 5'd0;
    frame0[28][14] = 5'd0;
    frame0[29][14] = 5'd0;
    frame0[30][14] = 5'd0;
    frame0[31][14] = 5'd0;
    frame0[0][15] = 5'd0;
    frame0[1][15] = 5'd0;
    frame0[2][15] = 5'd0;
    frame0[3][15] = 5'd0;
    frame0[4][15] = 5'd0;
    frame0[5][15] = 5'd0;
    frame0[6][15] = 5'd0;
    frame0[7][15] = 5'd0;
    frame0[8][15] = 5'd0;
    frame0[9][15] = 5'd0;
    frame0[10][15] = 5'd0;
    frame0[11][15] = 5'd0;
    frame0[12][15] = 5'd0;
    frame0[13][15] = 5'd0;
    frame0[14][15] = 5'd0;
    frame0[15][15] = 5'd0;
    frame0[16][15] = 5'd0;
    frame0[17][15] = 5'd0;
    frame0[18][15] = 5'd0;
    frame0[19][15] = 5'd0;
    frame0[20][15] = 5'd0;
    frame0[21][15] = 5'd0;
    frame0[22][15] = 5'd0;
    frame0[23][15] = 5'd0;
    frame0[24][15] = 5'd0;
    frame0[25][15] = 5'd0;
    frame0[26][15] = 5'd0;
    frame0[27][15] = 5'd0;
    frame0[28][15] = 5'd0;
    frame0[29][15] = 5'd0;
    frame0[30][15] = 5'd0;
    frame0[31][15] = 5'd0;
    frame0[0][16] = 5'd0;
    frame0[1][16] = 5'd0;
    frame0[2][16] = 5'd0;
    frame0[3][16] = 5'd0;
    frame0[4][16] = 5'd0;
    frame0[5][16] = 5'd0;
    frame0[6][16] = 5'd0;
    frame0[7][16] = 5'd0;
    frame0[8][16] = 5'd0;
    frame0[9][16] = 5'd0;
    frame0[10][16] = 5'd0;
    frame0[11][16] = 5'd0;
    frame0[12][16] = 5'd0;
    frame0[13][16] = 5'd0;
    frame0[14][16] = 5'd0;
    frame0[15][16] = 5'd0;
    frame0[16][16] = 5'd0;
    frame0[17][16] = 5'd0;
    frame0[18][16] = 5'd0;
    frame0[19][16] = 5'd0;
    frame0[20][16] = 5'd0;
    frame0[21][16] = 5'd0;
    frame0[22][16] = 5'd0;
    frame0[23][16] = 5'd0;
    frame0[24][16] = 5'd0;
    frame0[25][16] = 5'd0;
    frame0[26][16] = 5'd0;
    frame0[27][16] = 5'd0;
    frame0[28][16] = 5'd0;
    frame0[29][16] = 5'd0;
    frame0[30][16] = 5'd0;
    frame0[31][16] = 5'd0;
    frame0[0][17] = 5'd0;
    frame0[1][17] = 5'd0;
    frame0[2][17] = 5'd0;
    frame0[3][17] = 5'd0;
    frame0[4][17] = 5'd0;
    frame0[5][17] = 5'd0;
    frame0[6][17] = 5'd0;
    frame0[7][17] = 5'd0;
    frame0[8][17] = 5'd0;
    frame0[9][17] = 5'd0;
    frame0[10][17] = 5'd0;
    frame0[11][17] = 5'd0;
    frame0[12][17] = 5'd0;
    frame0[13][17] = 5'd0;
    frame0[14][17] = 5'd0;
    frame0[15][17] = 5'd0;
    frame0[16][17] = 5'd0;
    frame0[17][17] = 5'd0;
    frame0[18][17] = 5'd0;
    frame0[19][17] = 5'd0;
    frame0[20][17] = 5'd0;
    frame0[21][17] = 5'd0;
    frame0[22][17] = 5'd0;
    frame0[23][17] = 5'd0;
    frame0[24][17] = 5'd0;
    frame0[25][17] = 5'd0;
    frame0[26][17] = 5'd0;
    frame0[27][17] = 5'd0;
    frame0[28][17] = 5'd0;
    frame0[29][17] = 5'd0;
    frame0[30][17] = 5'd0;
    frame0[31][17] = 5'd0;
    frame0[0][18] = 5'd0;
    frame0[1][18] = 5'd0;
    frame0[2][18] = 5'd0;
    frame0[3][18] = 5'd0;
    frame0[4][18] = 5'd0;
    frame0[5][18] = 5'd0;
    frame0[6][18] = 5'd0;
    frame0[7][18] = 5'd0;
    frame0[8][18] = 5'd0;
    frame0[9][18] = 5'd0;
    frame0[10][18] = 5'd0;
    frame0[11][18] = 5'd0;
    frame0[12][18] = 5'd0;
    frame0[13][18] = 5'd0;
    frame0[14][18] = 5'd0;
    frame0[15][18] = 5'd0;
    frame0[16][18] = 5'd0;
    frame0[17][18] = 5'd0;
    frame0[18][18] = 5'd0;
    frame0[19][18] = 5'd0;
    frame0[20][18] = 5'd0;
    frame0[21][18] = 5'd0;
    frame0[22][18] = 5'd0;
    frame0[23][18] = 5'd0;
    frame0[24][18] = 5'd0;
    frame0[25][18] = 5'd0;
    frame0[26][18] = 5'd0;
    frame0[27][18] = 5'd0;
    frame0[28][18] = 5'd0;
    frame0[29][18] = 5'd0;
    frame0[30][18] = 5'd0;
    frame0[31][18] = 5'd0;
    frame0[0][19] = 5'd0;
    frame0[1][19] = 5'd0;
    frame0[2][19] = 5'd0;
    frame0[3][19] = 5'd0;
    frame0[4][19] = 5'd0;
    frame0[5][19] = 5'd0;
    frame0[6][19] = 5'd0;
    frame0[7][19] = 5'd0;
    frame0[8][19] = 5'd0;
    frame0[9][19] = 5'd0;
    frame0[10][19] = 5'd0;
    frame0[11][19] = 5'd0;
    frame0[12][19] = 5'd0;
    frame0[13][19] = 5'd0;
    frame0[14][19] = 5'd0;
    frame0[15][19] = 5'd0;
    frame0[16][19] = 5'd0;
    frame0[17][19] = 5'd0;
    frame0[18][19] = 5'd0;
    frame0[19][19] = 5'd0;
    frame0[20][19] = 5'd0;
    frame0[21][19] = 5'd0;
    frame0[22][19] = 5'd0;
    frame0[23][19] = 5'd0;
    frame0[24][19] = 5'd0;
    frame0[25][19] = 5'd0;
    frame0[26][19] = 5'd0;
    frame0[27][19] = 5'd0;
    frame0[28][19] = 5'd0;
    frame0[29][19] = 5'd0;
    frame0[30][19] = 5'd0;
    frame0[31][19] = 5'd0;
    frame0[0][20] = 5'd0;
    frame0[1][20] = 5'd0;
    frame0[2][20] = 5'd0;
    frame0[3][20] = 5'd0;
    frame0[4][20] = 5'd0;
    frame0[5][20] = 5'd0;
    frame0[6][20] = 5'd0;
    frame0[7][20] = 5'd0;
    frame0[8][20] = 5'd0;
    frame0[9][20] = 5'd0;
    frame0[10][20] = 5'd0;
    frame0[11][20] = 5'd0;
    frame0[12][20] = 5'd0;
    frame0[13][20] = 5'd0;
    frame0[14][20] = 5'd0;
    frame0[15][20] = 5'd0;
    frame0[16][20] = 5'd0;
    frame0[17][20] = 5'd0;
    frame0[18][20] = 5'd0;
    frame0[19][20] = 5'd0;
    frame0[20][20] = 5'd0;
    frame0[21][20] = 5'd0;
    frame0[22][20] = 5'd0;
    frame0[23][20] = 5'd0;
    frame0[24][20] = 5'd0;
    frame0[25][20] = 5'd0;
    frame0[26][20] = 5'd0;
    frame0[27][20] = 5'd0;
    frame0[28][20] = 5'd0;
    frame0[29][20] = 5'd0;
    frame0[30][20] = 5'd0;
    frame0[31][20] = 5'd0;
    frame0[0][21] = 5'd0;
    frame0[1][21] = 5'd0;
    frame0[2][21] = 5'd0;
    frame0[3][21] = 5'd0;
    frame0[4][21] = 5'd0;
    frame0[5][21] = 5'd0;
    frame0[6][21] = 5'd0;
    frame0[7][21] = 5'd0;
    frame0[8][21] = 5'd0;
    frame0[9][21] = 5'd0;
    frame0[10][21] = 5'd0;
    frame0[11][21] = 5'd0;
    frame0[12][21] = 5'd0;
    frame0[13][21] = 5'd0;
    frame0[14][21] = 5'd0;
    frame0[15][21] = 5'd0;
    frame0[16][21] = 5'd0;
    frame0[17][21] = 5'd0;
    frame0[18][21] = 5'd0;
    frame0[19][21] = 5'd0;
    frame0[20][21] = 5'd0;
    frame0[21][21] = 5'd0;
    frame0[22][21] = 5'd0;
    frame0[23][21] = 5'd0;
    frame0[24][21] = 5'd0;
    frame0[25][21] = 5'd0;
    frame0[26][21] = 5'd0;
    frame0[27][21] = 5'd0;
    frame0[28][21] = 5'd0;
    frame0[29][21] = 5'd0;
    frame0[30][21] = 5'd0;
    frame0[31][21] = 5'd0;
    frame0[0][22] = 5'd0;
    frame0[1][22] = 5'd0;
    frame0[2][22] = 5'd0;
    frame0[3][22] = 5'd0;
    frame0[4][22] = 5'd0;
    frame0[5][22] = 5'd0;
    frame0[6][22] = 5'd0;
    frame0[7][22] = 5'd0;
    frame0[8][22] = 5'd0;
    frame0[9][22] = 5'd0;
    frame0[10][22] = 5'd0;
    frame0[11][22] = 5'd0;
    frame0[12][22] = 5'd0;
    frame0[13][22] = 5'd0;
    frame0[14][22] = 5'd0;
    frame0[15][22] = 5'd0;
    frame0[16][22] = 5'd0;
    frame0[17][22] = 5'd0;
    frame0[18][22] = 5'd0;
    frame0[19][22] = 5'd0;
    frame0[20][22] = 5'd0;
    frame0[21][22] = 5'd0;
    frame0[22][22] = 5'd0;
    frame0[23][22] = 5'd0;
    frame0[24][22] = 5'd0;
    frame0[25][22] = 5'd0;
    frame0[26][22] = 5'd0;
    frame0[27][22] = 5'd0;
    frame0[28][22] = 5'd0;
    frame0[29][22] = 5'd0;
    frame0[30][22] = 5'd0;
    frame0[31][22] = 5'd0;
    frame0[0][23] = 5'd0;
    frame0[1][23] = 5'd0;
    frame0[2][23] = 5'd0;
    frame0[3][23] = 5'd0;
    frame0[4][23] = 5'd0;
    frame0[5][23] = 5'd0;
    frame0[6][23] = 5'd0;
    frame0[7][23] = 5'd0;
    frame0[8][23] = 5'd0;
    frame0[9][23] = 5'd0;
    frame0[10][23] = 5'd0;
    frame0[11][23] = 5'd0;
    frame0[12][23] = 5'd0;
    frame0[13][23] = 5'd0;
    frame0[14][23] = 5'd0;
    frame0[15][23] = 5'd0;
    frame0[16][23] = 5'd0;
    frame0[17][23] = 5'd0;
    frame0[18][23] = 5'd0;
    frame0[19][23] = 5'd0;
    frame0[20][23] = 5'd0;
    frame0[21][23] = 5'd0;
    frame0[22][23] = 5'd0;
    frame0[23][23] = 5'd0;
    frame0[24][23] = 5'd0;
    frame0[25][23] = 5'd0;
    frame0[26][23] = 5'd0;
    frame0[27][23] = 5'd0;
    frame0[28][23] = 5'd0;
    frame0[29][23] = 5'd0;
    frame0[30][23] = 5'd0;
    frame0[31][23] = 5'd0;
    frame0[0][24] = 5'd0;
    frame0[1][24] = 5'd0;
    frame0[2][24] = 5'd0;
    frame0[3][24] = 5'd0;
    frame0[4][24] = 5'd0;
    frame0[5][24] = 5'd0;
    frame0[6][24] = 5'd0;
    frame0[7][24] = 5'd0;
    frame0[8][24] = 5'd0;
    frame0[9][24] = 5'd0;
    frame0[10][24] = 5'd0;
    frame0[11][24] = 5'd0;
    frame0[12][24] = 5'd0;
    frame0[13][24] = 5'd0;
    frame0[14][24] = 5'd0;
    frame0[15][24] = 5'd0;
    frame0[16][24] = 5'd0;
    frame0[17][24] = 5'd0;
    frame0[18][24] = 5'd0;
    frame0[19][24] = 5'd0;
    frame0[20][24] = 5'd0;
    frame0[21][24] = 5'd0;
    frame0[22][24] = 5'd0;
    frame0[23][24] = 5'd0;
    frame0[24][24] = 5'd0;
    frame0[25][24] = 5'd0;
    frame0[26][24] = 5'd0;
    frame0[27][24] = 5'd0;
    frame0[28][24] = 5'd0;
    frame0[29][24] = 5'd0;
    frame0[30][24] = 5'd0;
    frame0[31][24] = 5'd0;
    frame0[0][25] = 5'd0;
    frame0[1][25] = 5'd0;
    frame0[2][25] = 5'd0;
    frame0[3][25] = 5'd0;
    frame0[4][25] = 5'd0;
    frame0[5][25] = 5'd0;
    frame0[6][25] = 5'd0;
    frame0[7][25] = 5'd0;
    frame0[8][25] = 5'd0;
    frame0[9][25] = 5'd0;
    frame0[10][25] = 5'd0;
    frame0[11][25] = 5'd0;
    frame0[12][25] = 5'd0;
    frame0[13][25] = 5'd0;
    frame0[14][25] = 5'd0;
    frame0[15][25] = 5'd0;
    frame0[16][25] = 5'd0;
    frame0[17][25] = 5'd0;
    frame0[18][25] = 5'd0;
    frame0[19][25] = 5'd0;
    frame0[20][25] = 5'd0;
    frame0[21][25] = 5'd0;
    frame0[22][25] = 5'd0;
    frame0[23][25] = 5'd0;
    frame0[24][25] = 5'd0;
    frame0[25][25] = 5'd0;
    frame0[26][25] = 5'd0;
    frame0[27][25] = 5'd0;
    frame0[28][25] = 5'd0;
    frame0[29][25] = 5'd0;
    frame0[30][25] = 5'd0;
    frame0[31][25] = 5'd0;
    frame0[0][26] = 5'd0;
    frame0[1][26] = 5'd0;
    frame0[2][26] = 5'd0;
    frame0[3][26] = 5'd0;
    frame0[4][26] = 5'd0;
    frame0[5][26] = 5'd0;
    frame0[6][26] = 5'd0;
    frame0[7][26] = 5'd0;
    frame0[8][26] = 5'd0;
    frame0[9][26] = 5'd0;
    frame0[10][26] = 5'd0;
    frame0[11][26] = 5'd0;
    frame0[12][26] = 5'd0;
    frame0[13][26] = 5'd0;
    frame0[14][26] = 5'd0;
    frame0[15][26] = 5'd0;
    frame0[16][26] = 5'd15;
    frame0[17][26] = 5'd3;
    frame0[18][26] = 5'd3;
    frame0[19][26] = 5'd3;
    frame0[20][26] = 5'd3;
    frame0[21][26] = 5'd3;
    frame0[22][26] = 5'd3;
    frame0[23][26] = 5'd3;
    frame0[24][26] = 5'd3;
    frame0[25][26] = 5'd0;
    frame0[26][26] = 5'd0;
    frame0[27][26] = 5'd0;
    frame0[28][26] = 5'd0;
    frame0[29][26] = 5'd0;
    frame0[30][26] = 5'd0;
    frame0[31][26] = 5'd0;
    frame0[0][27] = 5'd0;
    frame0[1][27] = 5'd0;
    frame0[2][27] = 5'd0;
    frame0[3][27] = 5'd0;
    frame0[4][27] = 5'd0;
    frame0[5][27] = 5'd0;
    frame0[6][27] = 5'd0;
    frame0[7][27] = 5'd0;
    frame0[8][27] = 5'd5;
    frame0[9][27] = 5'd5;
    frame0[10][27] = 5'd5;
    frame0[11][27] = 5'd5;
    frame0[12][27] = 5'd0;
    frame0[13][27] = 5'd0;
    frame0[14][27] = 5'd0;
    frame0[15][27] = 5'd0;
    frame0[16][27] = 5'd22;
    frame0[17][27] = 5'd9;
    frame0[18][27] = 5'd9;
    frame0[19][27] = 5'd9;
    frame0[20][27] = 5'd9;
    frame0[21][27] = 5'd9;
    frame0[22][27] = 5'd9;
    frame0[23][27] = 5'd9;
    frame0[24][27] = 5'd9;
    frame0[25][27] = 5'd14;
    frame0[26][27] = 5'd0;
    frame0[27][27] = 5'd0;
    frame0[28][27] = 5'd0;
    frame0[29][27] = 5'd0;
    frame0[30][27] = 5'd0;
    frame0[31][27] = 5'd0;
    frame0[0][28] = 5'd0;
    frame0[1][28] = 5'd0;
    frame0[2][28] = 5'd0;
    frame0[3][28] = 5'd0;
    frame0[4][28] = 5'd0;
    frame0[5][28] = 5'd0;
    frame0[6][28] = 5'd0;
    frame0[7][28] = 5'd0;
    frame0[8][28] = 5'd5;
    frame0[9][28] = 5'd5;
    frame0[10][28] = 5'd5;
    frame0[11][28] = 5'd5;
    frame0[12][28] = 5'd0;
    frame0[13][28] = 5'd0;
    frame0[14][28] = 5'd0;
    frame0[15][28] = 5'd15;
    frame0[16][28] = 5'd9;
    frame0[17][28] = 5'd13;
    frame0[18][28] = 5'd1;
    frame0[19][28] = 5'd1;
    frame0[20][28] = 5'd1;
    frame0[21][28] = 5'd1;
    frame0[22][28] = 5'd1;
    frame0[23][28] = 5'd1;
    frame0[24][28] = 5'd9;
    frame0[25][28] = 5'd16;
    frame0[26][28] = 5'd0;
    frame0[27][28] = 5'd0;
    frame0[28][28] = 5'd0;
    frame0[29][28] = 5'd0;
    frame0[30][28] = 5'd0;
    frame0[31][28] = 5'd0;
    frame0[0][29] = 5'd0;
    frame0[1][29] = 5'd0;
    frame0[2][29] = 5'd0;
    frame0[3][29] = 5'd0;
    frame0[4][29] = 5'd5;
    frame0[5][29] = 5'd5;
    frame0[6][29] = 5'd5;
    frame0[7][29] = 5'd5;
    frame0[8][29] = 5'd4;
    frame0[9][29] = 5'd4;
    frame0[10][29] = 5'd4;
    frame0[11][29] = 5'd4;
    frame0[12][29] = 5'd5;
    frame0[13][29] = 5'd5;
    frame0[14][29] = 5'd5;
    frame0[15][29] = 5'd21;
    frame0[16][29] = 5'd9;
    frame0[17][29] = 5'd1;
    frame0[18][29] = 5'd1;
    frame0[19][29] = 5'd1;
    frame0[20][29] = 5'd17;
    frame0[21][29] = 5'd19;
    frame0[22][29] = 5'd1;
    frame0[23][29] = 5'd1;
    frame0[24][29] = 5'd31;
    frame0[25][29] = 5'd16;
    frame0[26][29] = 5'd0;
    frame0[27][29] = 5'd0;
    frame0[28][29] = 5'd0;
    frame0[29][29] = 5'd0;
    frame0[30][29] = 5'd0;
    frame0[31][29] = 5'd0;
    frame0[0][30] = 5'd0;
    frame0[1][30] = 5'd0;
    frame0[2][30] = 5'd0;
    frame0[3][30] = 5'd0;
    frame0[4][30] = 5'd5;
    frame0[5][30] = 5'd5;
    frame0[6][30] = 5'd5;
    frame0[7][30] = 5'd5;
    frame0[8][30] = 5'd4;
    frame0[9][30] = 5'd4;
    frame0[10][30] = 5'd4;
    frame0[11][30] = 5'd4;
    frame0[12][30] = 5'd5;
    frame0[13][30] = 5'd5;
    frame0[14][30] = 5'd5;
    frame0[15][30] = 5'd21;
    frame0[16][30] = 5'd13;
    frame0[17][30] = 5'd19;
    frame0[18][30] = 5'd1;
    frame0[19][30] = 5'd1;
    frame0[20][30] = 5'd1;
    frame0[21][30] = 5'd1;
    frame0[22][30] = 5'd1;
    frame0[23][30] = 5'd1;
    frame0[24][30] = 5'd1;
    frame0[25][30] = 5'd16;
    frame0[26][30] = 5'd0;
    frame0[27][30] = 5'd0;
    frame0[28][30] = 5'd0;
    frame0[29][30] = 5'd0;
    frame0[30][30] = 5'd0;
    frame0[31][30] = 5'd0;
    frame0[0][31] = 5'd0;
    frame0[1][31] = 5'd0;
    frame0[2][31] = 5'd0;
    frame0[3][31] = 5'd0;
    frame0[4][31] = 5'd4;
    frame0[5][31] = 5'd4;
    frame0[6][31] = 5'd4;
    frame0[7][31] = 5'd4;
    frame0[8][31] = 5'd6;
    frame0[9][31] = 5'd6;
    frame0[10][31] = 5'd6;
    frame0[11][31] = 5'd6;
    frame0[12][31] = 5'd4;
    frame0[13][31] = 5'd4;
    frame0[14][31] = 5'd4;
    frame0[15][31] = 5'd28;
    frame0[16][31] = 5'd13;
    frame0[17][31] = 5'd1;
    frame0[18][31] = 5'd1;
    frame0[19][31] = 5'd1;
    frame0[20][31] = 5'd1;
    frame0[21][31] = 5'd1;
    frame0[22][31] = 5'd3;
    frame0[23][31] = 5'd19;
    frame0[24][31] = 5'd1;
    frame0[25][31] = 5'd16;
    frame0[26][31] = 5'd0;
    frame0[27][31] = 5'd3;
    frame0[28][31] = 5'd0;
    frame0[29][31] = 5'd0;
    frame0[30][31] = 5'd0;
    frame0[31][31] = 5'd0;
    frame0[0][32] = 5'd0;
    frame0[1][32] = 5'd0;
    frame0[2][32] = 5'd0;
    frame0[3][32] = 5'd0;
    frame0[4][32] = 5'd4;
    frame0[5][32] = 5'd4;
    frame0[6][32] = 5'd4;
    frame0[7][32] = 5'd4;
    frame0[8][32] = 5'd6;
    frame0[9][32] = 5'd6;
    frame0[10][32] = 5'd6;
    frame0[11][32] = 5'd6;
    frame0[12][32] = 5'd4;
    frame0[13][32] = 5'd4;
    frame0[14][32] = 5'd4;
    frame0[15][32] = 5'd28;
    frame0[16][32] = 5'd13;
    frame0[17][32] = 5'd1;
    frame0[18][32] = 5'd1;
    frame0[19][32] = 5'd1;
    frame0[20][32] = 5'd1;
    frame0[21][32] = 5'd18;
    frame0[22][32] = 5'd11;
    frame0[23][32] = 5'd1;
    frame0[24][32] = 5'd1;
    frame0[25][32] = 5'd16;
    frame0[26][32] = 5'd15;
    frame0[27][32] = 5'd2;
    frame0[28][32] = 5'd14;
    frame0[29][32] = 5'd0;
    frame0[30][32] = 5'd0;
    frame0[31][32] = 5'd0;
    frame0[0][33] = 5'd0;
    frame0[1][33] = 5'd0;
    frame0[2][33] = 5'd0;
    frame0[3][33] = 5'd0;
    frame0[4][33] = 5'd6;
    frame0[5][33] = 5'd6;
    frame0[6][33] = 5'd6;
    frame0[7][33] = 5'd6;
    frame0[8][33] = 5'd7;
    frame0[9][33] = 5'd7;
    frame0[10][33] = 5'd7;
    frame0[11][33] = 5'd7;
    frame0[12][33] = 5'd6;
    frame0[13][33] = 5'd6;
    frame0[14][33] = 5'd6;
    frame0[15][33] = 5'd23;
    frame0[16][33] = 5'd13;
    frame0[17][33] = 5'd1;
    frame0[18][33] = 5'd1;
    frame0[19][33] = 5'd19;
    frame0[20][33] = 5'd1;
    frame0[21][33] = 5'd18;
    frame0[22][33] = 5'd2;
    frame0[23][33] = 5'd3;
    frame0[24][33] = 5'd1;
    frame0[25][33] = 5'd16;
    frame0[26][33] = 5'd12;
    frame0[27][33] = 5'd2;
    frame0[28][33] = 5'd14;
    frame0[29][33] = 5'd0;
    frame0[30][33] = 5'd0;
    frame0[31][33] = 5'd0;
    frame0[0][34] = 5'd0;
    frame0[1][34] = 5'd0;
    frame0[2][34] = 5'd0;
    frame0[3][34] = 5'd0;
    frame0[4][34] = 5'd6;
    frame0[5][34] = 5'd6;
    frame0[6][34] = 5'd6;
    frame0[7][34] = 5'd6;
    frame0[8][34] = 5'd7;
    frame0[9][34] = 5'd7;
    frame0[10][34] = 5'd7;
    frame0[11][34] = 5'd7;
    frame0[12][34] = 5'd6;
    frame0[13][34] = 5'd3;
    frame0[14][34] = 5'd6;
    frame0[15][34] = 5'd23;
    frame0[16][34] = 5'd13;
    frame0[17][34] = 5'd1;
    frame0[18][34] = 5'd1;
    frame0[19][34] = 5'd1;
    frame0[20][34] = 5'd1;
    frame0[21][34] = 5'd18;
    frame0[22][34] = 5'd2;
    frame0[23][34] = 5'd2;
    frame0[24][34] = 5'd3;
    frame0[25][34] = 5'd3;
    frame0[26][34] = 5'd2;
    frame0[27][34] = 5'd2;
    frame0[28][34] = 5'd14;
    frame0[29][34] = 5'd0;
    frame0[30][34] = 5'd0;
    frame0[31][34] = 5'd0;
    frame0[0][35] = 5'd0;
    frame0[1][35] = 5'd0;
    frame0[2][35] = 5'd0;
    frame0[3][35] = 5'd0;
    frame0[4][35] = 5'd7;
    frame0[5][35] = 5'd7;
    frame0[6][35] = 5'd7;
    frame0[7][35] = 5'd7;
    frame0[8][35] = 5'd10;
    frame0[9][35] = 5'd10;
    frame0[10][35] = 5'd10;
    frame0[11][35] = 5'd10;
    frame0[12][35] = 5'd24;
    frame0[13][35] = 5'd11;
    frame0[14][35] = 5'd7;
    frame0[15][35] = 5'd24;
    frame0[16][35] = 5'd13;
    frame0[17][35] = 5'd1;
    frame0[18][35] = 5'd17;
    frame0[19][35] = 5'd1;
    frame0[20][35] = 5'd1;
    frame0[21][35] = 5'd18;
    frame0[22][35] = 5'd2;
    frame0[23][35] = 5'd2;
    frame0[24][35] = 5'd2;
    frame0[25][35] = 5'd2;
    frame0[26][35] = 5'd2;
    frame0[27][35] = 5'd2;
    frame0[28][35] = 5'd14;
    frame0[29][35] = 5'd0;
    frame0[30][35] = 5'd0;
    frame0[31][35] = 5'd0;
    frame0[0][36] = 5'd0;
    frame0[1][36] = 5'd0;
    frame0[2][36] = 5'd0;
    frame0[3][36] = 5'd0;
    frame0[4][36] = 5'd7;
    frame0[5][36] = 5'd7;
    frame0[6][36] = 5'd7;
    frame0[7][36] = 5'd7;
    frame0[8][36] = 5'd10;
    frame0[9][36] = 5'd10;
    frame0[10][36] = 5'd10;
    frame0[11][36] = 5'd10;
    frame0[12][36] = 5'd24;
    frame0[13][36] = 5'd2;
    frame0[14][36] = 5'd3;
    frame0[15][36] = 5'd3;
    frame0[16][36] = 5'd13;
    frame0[17][36] = 5'd1;
    frame0[18][36] = 5'd1;
    frame0[19][36] = 5'd1;
    frame0[20][36] = 5'd17;
    frame0[21][36] = 5'd12;
    frame0[22][36] = 5'd2;
    frame0[23][36] = 5'd2;
    frame0[24][36] = 5'd2;
    frame0[25][36] = 5'd2;
    frame0[26][36] = 5'd2;
    frame0[27][36] = 5'd2;
    frame0[28][36] = 5'd11;
    frame0[29][36] = 5'd0;
    frame0[30][36] = 5'd0;
    frame0[31][36] = 5'd0;
    frame0[0][37] = 5'd0;
    frame0[1][37] = 5'd0;
    frame0[2][37] = 5'd0;
    frame0[3][37] = 5'd0;
    frame0[4][37] = 5'd10;
    frame0[5][37] = 5'd10;
    frame0[6][37] = 5'd10;
    frame0[7][37] = 5'd10;
    frame0[8][37] = 5'd8;
    frame0[9][37] = 5'd8;
    frame0[10][37] = 5'd8;
    frame0[11][37] = 5'd8;
    frame0[12][37] = 5'd10;
    frame0[13][37] = 5'd12;
    frame0[14][37] = 5'd2;
    frame0[15][37] = 5'd11;
    frame0[16][37] = 5'd13;
    frame0[17][37] = 5'd17;
    frame0[18][37] = 5'd1;
    frame0[19][37] = 5'd1;
    frame0[20][37] = 5'd1;
    frame0[21][37] = 5'd12;
    frame0[22][37] = 5'd2;
    frame0[23][37] = 5'd20;
    frame0[24][37] = 5'd2;
    frame0[25][37] = 5'd2;
    frame0[26][37] = 5'd20;
    frame0[27][37] = 5'd2;
    frame0[28][37] = 5'd11;
    frame0[29][37] = 5'd0;
    frame0[30][37] = 5'd0;
    frame0[31][37] = 5'd0;
    frame0[0][38] = 5'd0;
    frame0[1][38] = 5'd0;
    frame0[2][38] = 5'd0;
    frame0[3][38] = 5'd0;
    frame0[4][38] = 5'd10;
    frame0[5][38] = 5'd10;
    frame0[6][38] = 5'd10;
    frame0[7][38] = 5'd10;
    frame0[8][38] = 5'd8;
    frame0[9][38] = 5'd8;
    frame0[10][38] = 5'd8;
    frame0[11][38] = 5'd8;
    frame0[12][38] = 5'd10;
    frame0[13][38] = 5'd30;
    frame0[14][38] = 5'd12;
    frame0[15][38] = 5'd11;
    frame0[16][38] = 5'd13;
    frame0[17][38] = 5'd1;
    frame0[18][38] = 5'd1;
    frame0[19][38] = 5'd1;
    frame0[20][38] = 5'd1;
    frame0[21][38] = 5'd12;
    frame0[22][38] = 5'd2;
    frame0[23][38] = 5'd3;
    frame0[24][38] = 5'd2;
    frame0[25][38] = 5'd12;
    frame0[26][38] = 5'd3;
    frame0[27][38] = 5'd2;
    frame0[28][38] = 5'd11;
    frame0[29][38] = 5'd0;
    frame0[30][38] = 5'd0;
    frame0[31][38] = 5'd0;
    frame0[0][39] = 5'd0;
    frame0[1][39] = 5'd0;
    frame0[2][39] = 5'd0;
    frame0[3][39] = 5'd0;
    frame0[4][39] = 5'd8;
    frame0[5][39] = 5'd8;
    frame0[6][39] = 5'd8;
    frame0[7][39] = 5'd8;
    frame0[8][39] = 5'd0;
    frame0[9][39] = 5'd0;
    frame0[10][39] = 5'd0;
    frame0[11][39] = 5'd0;
    frame0[12][39] = 5'd8;
    frame0[13][39] = 5'd8;
    frame0[14][39] = 5'd29;
    frame0[15][39] = 5'd3;
    frame0[16][39] = 5'd13;
    frame0[17][39] = 5'd1;
    frame0[18][39] = 5'd1;
    frame0[19][39] = 5'd17;
    frame0[20][39] = 5'd1;
    frame0[21][39] = 5'd12;
    frame0[22][39] = 5'd25;
    frame0[23][39] = 5'd2;
    frame0[24][39] = 5'd2;
    frame0[25][39] = 5'd2;
    frame0[26][39] = 5'd2;
    frame0[27][39] = 5'd27;
    frame0[28][39] = 5'd26;
    frame0[29][39] = 5'd0;
    frame0[30][39] = 5'd0;
    frame0[31][39] = 5'd0;
    frame0[0][40] = 5'd0;
    frame0[1][40] = 5'd0;
    frame0[2][40] = 5'd0;
    frame0[3][40] = 5'd0;
    frame0[4][40] = 5'd8;
    frame0[5][40] = 5'd8;
    frame0[6][40] = 5'd8;
    frame0[7][40] = 5'd8;
    frame0[8][40] = 5'd0;
    frame0[9][40] = 5'd0;
    frame0[10][40] = 5'd0;
    frame0[11][40] = 5'd0;
    frame0[12][40] = 5'd8;
    frame0[13][40] = 5'd8;
    frame0[14][40] = 5'd8;
    frame0[15][40] = 5'd29;
    frame0[16][40] = 5'd9;
    frame0[17][40] = 5'd19;
    frame0[18][40] = 5'd1;
    frame0[19][40] = 5'd1;
    frame0[20][40] = 5'd1;
    frame0[21][40] = 5'd12;
    frame0[22][40] = 5'd25;
    frame0[23][40] = 5'd11;
    frame0[24][40] = 5'd2;
    frame0[25][40] = 5'd12;
    frame0[26][40] = 5'd11;
    frame0[27][40] = 5'd27;
    frame0[28][40] = 5'd26;
    frame0[29][40] = 5'd0;
    frame0[30][40] = 5'd0;
    frame0[31][40] = 5'd0;
    frame0[0][41] = 5'd0;
    frame0[1][41] = 5'd0;
    frame0[2][41] = 5'd0;
    frame0[3][41] = 5'd0;
    frame0[4][41] = 5'd0;
    frame0[5][41] = 5'd0;
    frame0[6][41] = 5'd0;
    frame0[7][41] = 5'd0;
    frame0[8][41] = 5'd0;
    frame0[9][41] = 5'd0;
    frame0[10][41] = 5'd0;
    frame0[11][41] = 5'd0;
    frame0[12][41] = 5'd0;
    frame0[13][41] = 5'd0;
    frame0[14][41] = 5'd0;
    frame0[15][41] = 5'd15;
    frame0[16][41] = 5'd9;
    frame0[17][41] = 5'd13;
    frame0[18][41] = 5'd1;
    frame0[19][41] = 5'd1;
    frame0[20][41] = 5'd1;
    frame0[21][41] = 5'd18;
    frame0[22][41] = 5'd2;
    frame0[23][41] = 5'd11;
    frame0[24][41] = 5'd3;
    frame0[25][41] = 5'd3;
    frame0[26][41] = 5'd3;
    frame0[27][41] = 5'd2;
    frame0[28][41] = 5'd14;
    frame0[29][41] = 5'd0;
    frame0[30][41] = 5'd0;
    frame0[31][41] = 5'd0;
    frame0[0][42] = 5'd0;
    frame0[1][42] = 5'd0;
    frame0[2][42] = 5'd0;
    frame0[3][42] = 5'd0;
    frame0[4][42] = 5'd0;
    frame0[5][42] = 5'd0;
    frame0[6][42] = 5'd0;
    frame0[7][42] = 5'd0;
    frame0[8][42] = 5'd0;
    frame0[9][42] = 5'd0;
    frame0[10][42] = 5'd0;
    frame0[11][42] = 5'd0;
    frame0[12][42] = 5'd0;
    frame0[13][42] = 5'd0;
    frame0[14][42] = 5'd0;
    frame0[15][42] = 5'd15;
    frame0[16][42] = 5'd22;
    frame0[17][42] = 5'd9;
    frame0[18][42] = 5'd9;
    frame0[19][42] = 5'd9;
    frame0[20][42] = 5'd9;
    frame0[21][42] = 5'd9;
    frame0[22][42] = 5'd12;
    frame0[23][42] = 5'd2;
    frame0[24][42] = 5'd2;
    frame0[25][42] = 5'd2;
    frame0[26][42] = 5'd2;
    frame0[27][42] = 5'd11;
    frame0[28][42] = 5'd0;
    frame0[29][42] = 5'd0;
    frame0[30][42] = 5'd0;
    frame0[31][42] = 5'd0;
    frame0[0][43] = 5'd0;
    frame0[1][43] = 5'd0;
    frame0[2][43] = 5'd0;
    frame0[3][43] = 5'd0;
    frame0[4][43] = 5'd0;
    frame0[5][43] = 5'd0;
    frame0[6][43] = 5'd0;
    frame0[7][43] = 5'd0;
    frame0[8][43] = 5'd0;
    frame0[9][43] = 5'd0;
    frame0[10][43] = 5'd0;
    frame0[11][43] = 5'd0;
    frame0[12][43] = 5'd0;
    frame0[13][43] = 5'd0;
    frame0[14][43] = 5'd0;
    frame0[15][43] = 5'd15;
    frame0[16][43] = 5'd11;
    frame0[17][43] = 5'd3;
    frame0[18][43] = 5'd3;
    frame0[19][43] = 5'd3;
    frame0[20][43] = 5'd3;
    frame0[21][43] = 5'd3;
    frame0[22][43] = 5'd3;
    frame0[23][43] = 5'd3;
    frame0[24][43] = 5'd3;
    frame0[25][43] = 5'd3;
    frame0[26][43] = 5'd3;
    frame0[27][43] = 5'd14;
    frame0[28][43] = 5'd0;
    frame0[29][43] = 5'd0;
    frame0[30][43] = 5'd0;
    frame0[31][43] = 5'd0;
    frame0[0][44] = 5'd0;
    frame0[1][44] = 5'd0;
    frame0[2][44] = 5'd0;
    frame0[3][44] = 5'd0;
    frame0[4][44] = 5'd0;
    frame0[5][44] = 5'd0;
    frame0[6][44] = 5'd0;
    frame0[7][44] = 5'd0;
    frame0[8][44] = 5'd0;
    frame0[9][44] = 5'd0;
    frame0[10][44] = 5'd0;
    frame0[11][44] = 5'd0;
    frame0[12][44] = 5'd0;
    frame0[13][44] = 5'd0;
    frame0[14][44] = 5'd0;
    frame0[15][44] = 5'd15;
    frame0[16][44] = 5'd2;
    frame0[17][44] = 5'd14;
    frame0[18][44] = 5'd12;
    frame0[19][44] = 5'd11;
    frame0[20][44] = 5'd0;
    frame0[21][44] = 5'd0;
    frame0[22][44] = 5'd0;
    frame0[23][44] = 5'd12;
    frame0[24][44] = 5'd11;
    frame0[25][44] = 5'd15;
    frame0[26][44] = 5'd2;
    frame0[27][44] = 5'd14;
    frame0[28][44] = 5'd0;
    frame0[29][44] = 5'd0;
    frame0[30][44] = 5'd0;
    frame0[31][44] = 5'd0;
    frame0[0][45] = 5'd0;
    frame0[1][45] = 5'd0;
    frame0[2][45] = 5'd0;
    frame0[3][45] = 5'd0;
    frame0[4][45] = 5'd0;
    frame0[5][45] = 5'd0;
    frame0[6][45] = 5'd0;
    frame0[7][45] = 5'd0;
    frame0[8][45] = 5'd0;
    frame0[9][45] = 5'd0;
    frame0[10][45] = 5'd0;
    frame0[11][45] = 5'd0;
    frame0[12][45] = 5'd0;
    frame0[13][45] = 5'd0;
    frame0[14][45] = 5'd0;
    frame0[15][45] = 5'd15;
    frame0[16][45] = 5'd3;
    frame0[17][45] = 5'd0;
    frame0[18][45] = 5'd15;
    frame0[19][45] = 5'd3;
    frame0[20][45] = 5'd0;
    frame0[21][45] = 5'd0;
    frame0[22][45] = 5'd0;
    frame0[23][45] = 5'd15;
    frame0[24][45] = 5'd3;
    frame0[25][45] = 5'd0;
    frame0[26][45] = 5'd3;
    frame0[27][45] = 5'd14;
    frame0[28][45] = 5'd0;
    frame0[29][45] = 5'd0;
    frame0[30][45] = 5'd0;
    frame0[31][45] = 5'd0;
    frame0[0][46] = 5'd0;
    frame0[1][46] = 5'd0;
    frame0[2][46] = 5'd0;
    frame0[3][46] = 5'd0;
    frame0[4][46] = 5'd0;
    frame0[5][46] = 5'd0;
    frame0[6][46] = 5'd0;
    frame0[7][46] = 5'd0;
    frame0[8][46] = 5'd0;
    frame0[9][46] = 5'd0;
    frame0[10][46] = 5'd0;
    frame0[11][46] = 5'd0;
    frame0[12][46] = 5'd0;
    frame0[13][46] = 5'd0;
    frame0[14][46] = 5'd0;
    frame0[15][46] = 5'd0;
    frame0[16][46] = 5'd0;
    frame0[17][46] = 5'd0;
    frame0[18][46] = 5'd0;
    frame0[19][46] = 5'd0;
    frame0[20][46] = 5'd0;
    frame0[21][46] = 5'd0;
    frame0[22][46] = 5'd0;
    frame0[23][46] = 5'd0;
    frame0[24][46] = 5'd0;
    frame0[25][46] = 5'd0;
    frame0[26][46] = 5'd0;
    frame0[27][46] = 5'd0;
    frame0[28][46] = 5'd0;
    frame0[29][46] = 5'd0;
    frame0[30][46] = 5'd0;
    frame0[31][46] = 5'd0;
    frame0[0][47] = 5'd0;
    frame0[1][47] = 5'd0;
    frame0[2][47] = 5'd0;
    frame0[3][47] = 5'd0;
    frame0[4][47] = 5'd0;
    frame0[5][47] = 5'd0;
    frame0[6][47] = 5'd0;
    frame0[7][47] = 5'd0;
    frame0[8][47] = 5'd0;
    frame0[9][47] = 5'd0;
    frame0[10][47] = 5'd0;
    frame0[11][47] = 5'd0;
    frame0[12][47] = 5'd0;
    frame0[13][47] = 5'd0;
    frame0[14][47] = 5'd0;
    frame0[15][47] = 5'd0;
    frame0[16][47] = 5'd0;
    frame0[17][47] = 5'd0;
    frame0[18][47] = 5'd0;
    frame0[19][47] = 5'd0;
    frame0[20][47] = 5'd0;
    frame0[21][47] = 5'd0;
    frame0[22][47] = 5'd0;
    frame0[23][47] = 5'd0;
    frame0[24][47] = 5'd0;
    frame0[25][47] = 5'd0;
    frame0[26][47] = 5'd0;
    frame0[27][47] = 5'd0;
    frame0[28][47] = 5'd0;
    frame0[29][47] = 5'd0;
    frame0[30][47] = 5'd0;
    frame0[31][47] = 5'd0;
end

reg [4:0] frame1[31:0][47:0];
initial begin
    frame1[0][0] = 5'd0;
    frame1[1][0] = 5'd0;
    frame1[2][0] = 5'd0;
    frame1[3][0] = 5'd0;
    frame1[4][0] = 5'd0;
    frame1[5][0] = 5'd0;
    frame1[6][0] = 5'd0;
    frame1[7][0] = 5'd0;
    frame1[8][0] = 5'd0;
    frame1[9][0] = 5'd0;
    frame1[10][0] = 5'd0;
    frame1[11][0] = 5'd0;
    frame1[12][0] = 5'd0;
    frame1[13][0] = 5'd0;
    frame1[14][0] = 5'd0;
    frame1[15][0] = 5'd0;
    frame1[16][0] = 5'd0;
    frame1[17][0] = 5'd0;
    frame1[18][0] = 5'd0;
    frame1[19][0] = 5'd0;
    frame1[20][0] = 5'd0;
    frame1[21][0] = 5'd0;
    frame1[22][0] = 5'd0;
    frame1[23][0] = 5'd0;
    frame1[24][0] = 5'd0;
    frame1[25][0] = 5'd0;
    frame1[26][0] = 5'd0;
    frame1[27][0] = 5'd0;
    frame1[28][0] = 5'd0;
    frame1[29][0] = 5'd0;
    frame1[30][0] = 5'd0;
    frame1[31][0] = 5'd0;
    frame1[0][1] = 5'd0;
    frame1[1][1] = 5'd0;
    frame1[2][1] = 5'd0;
    frame1[3][1] = 5'd0;
    frame1[4][1] = 5'd0;
    frame1[5][1] = 5'd0;
    frame1[6][1] = 5'd0;
    frame1[7][1] = 5'd0;
    frame1[8][1] = 5'd0;
    frame1[9][1] = 5'd0;
    frame1[10][1] = 5'd0;
    frame1[11][1] = 5'd0;
    frame1[12][1] = 5'd0;
    frame1[13][1] = 5'd0;
    frame1[14][1] = 5'd0;
    frame1[15][1] = 5'd0;
    frame1[16][1] = 5'd0;
    frame1[17][1] = 5'd0;
    frame1[18][1] = 5'd0;
    frame1[19][1] = 5'd0;
    frame1[20][1] = 5'd0;
    frame1[21][1] = 5'd0;
    frame1[22][1] = 5'd0;
    frame1[23][1] = 5'd0;
    frame1[24][1] = 5'd0;
    frame1[25][1] = 5'd0;
    frame1[26][1] = 5'd0;
    frame1[27][1] = 5'd0;
    frame1[28][1] = 5'd0;
    frame1[29][1] = 5'd0;
    frame1[30][1] = 5'd0;
    frame1[31][1] = 5'd0;
    frame1[0][2] = 5'd0;
    frame1[1][2] = 5'd0;
    frame1[2][2] = 5'd0;
    frame1[3][2] = 5'd0;
    frame1[4][2] = 5'd0;
    frame1[5][2] = 5'd0;
    frame1[6][2] = 5'd0;
    frame1[7][2] = 5'd0;
    frame1[8][2] = 5'd0;
    frame1[9][2] = 5'd0;
    frame1[10][2] = 5'd0;
    frame1[11][2] = 5'd0;
    frame1[12][2] = 5'd0;
    frame1[13][2] = 5'd0;
    frame1[14][2] = 5'd0;
    frame1[15][2] = 5'd0;
    frame1[16][2] = 5'd0;
    frame1[17][2] = 5'd0;
    frame1[18][2] = 5'd0;
    frame1[19][2] = 5'd0;
    frame1[20][2] = 5'd0;
    frame1[21][2] = 5'd0;
    frame1[22][2] = 5'd0;
    frame1[23][2] = 5'd0;
    frame1[24][2] = 5'd0;
    frame1[25][2] = 5'd0;
    frame1[26][2] = 5'd0;
    frame1[27][2] = 5'd0;
    frame1[28][2] = 5'd0;
    frame1[29][2] = 5'd0;
    frame1[30][2] = 5'd0;
    frame1[31][2] = 5'd0;
    frame1[0][3] = 5'd0;
    frame1[1][3] = 5'd0;
    frame1[2][3] = 5'd0;
    frame1[3][3] = 5'd0;
    frame1[4][3] = 5'd0;
    frame1[5][3] = 5'd0;
    frame1[6][3] = 5'd0;
    frame1[7][3] = 5'd0;
    frame1[8][3] = 5'd0;
    frame1[9][3] = 5'd0;
    frame1[10][3] = 5'd0;
    frame1[11][3] = 5'd0;
    frame1[12][3] = 5'd0;
    frame1[13][3] = 5'd0;
    frame1[14][3] = 5'd0;
    frame1[15][3] = 5'd0;
    frame1[16][3] = 5'd0;
    frame1[17][3] = 5'd0;
    frame1[18][3] = 5'd0;
    frame1[19][3] = 5'd0;
    frame1[20][3] = 5'd0;
    frame1[21][3] = 5'd0;
    frame1[22][3] = 5'd0;
    frame1[23][3] = 5'd0;
    frame1[24][3] = 5'd0;
    frame1[25][3] = 5'd0;
    frame1[26][3] = 5'd0;
    frame1[27][3] = 5'd0;
    frame1[28][3] = 5'd0;
    frame1[29][3] = 5'd0;
    frame1[30][3] = 5'd0;
    frame1[31][3] = 5'd0;
    frame1[0][4] = 5'd0;
    frame1[1][4] = 5'd0;
    frame1[2][4] = 5'd0;
    frame1[3][4] = 5'd0;
    frame1[4][4] = 5'd0;
    frame1[5][4] = 5'd0;
    frame1[6][4] = 5'd0;
    frame1[7][4] = 5'd0;
    frame1[8][4] = 5'd0;
    frame1[9][4] = 5'd0;
    frame1[10][4] = 5'd0;
    frame1[11][4] = 5'd0;
    frame1[12][4] = 5'd0;
    frame1[13][4] = 5'd0;
    frame1[14][4] = 5'd0;
    frame1[15][4] = 5'd0;
    frame1[16][4] = 5'd0;
    frame1[17][4] = 5'd0;
    frame1[18][4] = 5'd0;
    frame1[19][4] = 5'd0;
    frame1[20][4] = 5'd0;
    frame1[21][4] = 5'd0;
    frame1[22][4] = 5'd0;
    frame1[23][4] = 5'd0;
    frame1[24][4] = 5'd0;
    frame1[25][4] = 5'd0;
    frame1[26][4] = 5'd0;
    frame1[27][4] = 5'd0;
    frame1[28][4] = 5'd0;
    frame1[29][4] = 5'd0;
    frame1[30][4] = 5'd0;
    frame1[31][4] = 5'd0;
    frame1[0][5] = 5'd0;
    frame1[1][5] = 5'd0;
    frame1[2][5] = 5'd0;
    frame1[3][5] = 5'd0;
    frame1[4][5] = 5'd0;
    frame1[5][5] = 5'd0;
    frame1[6][5] = 5'd0;
    frame1[7][5] = 5'd0;
    frame1[8][5] = 5'd0;
    frame1[9][5] = 5'd0;
    frame1[10][5] = 5'd0;
    frame1[11][5] = 5'd0;
    frame1[12][5] = 5'd0;
    frame1[13][5] = 5'd0;
    frame1[14][5] = 5'd0;
    frame1[15][5] = 5'd0;
    frame1[16][5] = 5'd0;
    frame1[17][5] = 5'd0;
    frame1[18][5] = 5'd0;
    frame1[19][5] = 5'd0;
    frame1[20][5] = 5'd0;
    frame1[21][5] = 5'd0;
    frame1[22][5] = 5'd0;
    frame1[23][5] = 5'd0;
    frame1[24][5] = 5'd0;
    frame1[25][5] = 5'd0;
    frame1[26][5] = 5'd0;
    frame1[27][5] = 5'd0;
    frame1[28][5] = 5'd0;
    frame1[29][5] = 5'd0;
    frame1[30][5] = 5'd0;
    frame1[31][5] = 5'd0;
    frame1[0][6] = 5'd0;
    frame1[1][6] = 5'd0;
    frame1[2][6] = 5'd0;
    frame1[3][6] = 5'd0;
    frame1[4][6] = 5'd0;
    frame1[5][6] = 5'd0;
    frame1[6][6] = 5'd0;
    frame1[7][6] = 5'd0;
    frame1[8][6] = 5'd0;
    frame1[9][6] = 5'd0;
    frame1[10][6] = 5'd0;
    frame1[11][6] = 5'd0;
    frame1[12][6] = 5'd0;
    frame1[13][6] = 5'd0;
    frame1[14][6] = 5'd0;
    frame1[15][6] = 5'd0;
    frame1[16][6] = 5'd0;
    frame1[17][6] = 5'd0;
    frame1[18][6] = 5'd0;
    frame1[19][6] = 5'd0;
    frame1[20][6] = 5'd0;
    frame1[21][6] = 5'd0;
    frame1[22][6] = 5'd0;
    frame1[23][6] = 5'd0;
    frame1[24][6] = 5'd0;
    frame1[25][6] = 5'd0;
    frame1[26][6] = 5'd0;
    frame1[27][6] = 5'd0;
    frame1[28][6] = 5'd0;
    frame1[29][6] = 5'd0;
    frame1[30][6] = 5'd0;
    frame1[31][6] = 5'd0;
    frame1[0][7] = 5'd0;
    frame1[1][7] = 5'd0;
    frame1[2][7] = 5'd0;
    frame1[3][7] = 5'd0;
    frame1[4][7] = 5'd0;
    frame1[5][7] = 5'd0;
    frame1[6][7] = 5'd0;
    frame1[7][7] = 5'd0;
    frame1[8][7] = 5'd0;
    frame1[9][7] = 5'd0;
    frame1[10][7] = 5'd0;
    frame1[11][7] = 5'd0;
    frame1[12][7] = 5'd0;
    frame1[13][7] = 5'd0;
    frame1[14][7] = 5'd0;
    frame1[15][7] = 5'd0;
    frame1[16][7] = 5'd0;
    frame1[17][7] = 5'd0;
    frame1[18][7] = 5'd0;
    frame1[19][7] = 5'd0;
    frame1[20][7] = 5'd0;
    frame1[21][7] = 5'd0;
    frame1[22][7] = 5'd0;
    frame1[23][7] = 5'd0;
    frame1[24][7] = 5'd0;
    frame1[25][7] = 5'd0;
    frame1[26][7] = 5'd0;
    frame1[27][7] = 5'd0;
    frame1[28][7] = 5'd0;
    frame1[29][7] = 5'd0;
    frame1[30][7] = 5'd0;
    frame1[31][7] = 5'd0;
    frame1[0][8] = 5'd0;
    frame1[1][8] = 5'd0;
    frame1[2][8] = 5'd0;
    frame1[3][8] = 5'd0;
    frame1[4][8] = 5'd0;
    frame1[5][8] = 5'd0;
    frame1[6][8] = 5'd0;
    frame1[7][8] = 5'd0;
    frame1[8][8] = 5'd0;
    frame1[9][8] = 5'd0;
    frame1[10][8] = 5'd0;
    frame1[11][8] = 5'd0;
    frame1[12][8] = 5'd0;
    frame1[13][8] = 5'd0;
    frame1[14][8] = 5'd0;
    frame1[15][8] = 5'd0;
    frame1[16][8] = 5'd0;
    frame1[17][8] = 5'd0;
    frame1[18][8] = 5'd0;
    frame1[19][8] = 5'd0;
    frame1[20][8] = 5'd0;
    frame1[21][8] = 5'd0;
    frame1[22][8] = 5'd0;
    frame1[23][8] = 5'd0;
    frame1[24][8] = 5'd0;
    frame1[25][8] = 5'd0;
    frame1[26][8] = 5'd0;
    frame1[27][8] = 5'd0;
    frame1[28][8] = 5'd0;
    frame1[29][8] = 5'd0;
    frame1[30][8] = 5'd0;
    frame1[31][8] = 5'd0;
    frame1[0][9] = 5'd0;
    frame1[1][9] = 5'd0;
    frame1[2][9] = 5'd0;
    frame1[3][9] = 5'd0;
    frame1[4][9] = 5'd0;
    frame1[5][9] = 5'd0;
    frame1[6][9] = 5'd0;
    frame1[7][9] = 5'd0;
    frame1[8][9] = 5'd0;
    frame1[9][9] = 5'd0;
    frame1[10][9] = 5'd0;
    frame1[11][9] = 5'd0;
    frame1[12][9] = 5'd0;
    frame1[13][9] = 5'd0;
    frame1[14][9] = 5'd0;
    frame1[15][9] = 5'd0;
    frame1[16][9] = 5'd0;
    frame1[17][9] = 5'd0;
    frame1[18][9] = 5'd0;
    frame1[19][9] = 5'd0;
    frame1[20][9] = 5'd0;
    frame1[21][9] = 5'd0;
    frame1[22][9] = 5'd0;
    frame1[23][9] = 5'd0;
    frame1[24][9] = 5'd0;
    frame1[25][9] = 5'd0;
    frame1[26][9] = 5'd0;
    frame1[27][9] = 5'd0;
    frame1[28][9] = 5'd0;
    frame1[29][9] = 5'd0;
    frame1[30][9] = 5'd0;
    frame1[31][9] = 5'd0;
    frame1[0][10] = 5'd0;
    frame1[1][10] = 5'd0;
    frame1[2][10] = 5'd0;
    frame1[3][10] = 5'd0;
    frame1[4][10] = 5'd0;
    frame1[5][10] = 5'd0;
    frame1[6][10] = 5'd0;
    frame1[7][10] = 5'd0;
    frame1[8][10] = 5'd0;
    frame1[9][10] = 5'd0;
    frame1[10][10] = 5'd0;
    frame1[11][10] = 5'd0;
    frame1[12][10] = 5'd0;
    frame1[13][10] = 5'd0;
    frame1[14][10] = 5'd0;
    frame1[15][10] = 5'd0;
    frame1[16][10] = 5'd0;
    frame1[17][10] = 5'd0;
    frame1[18][10] = 5'd0;
    frame1[19][10] = 5'd0;
    frame1[20][10] = 5'd0;
    frame1[21][10] = 5'd0;
    frame1[22][10] = 5'd0;
    frame1[23][10] = 5'd0;
    frame1[24][10] = 5'd0;
    frame1[25][10] = 5'd0;
    frame1[26][10] = 5'd0;
    frame1[27][10] = 5'd0;
    frame1[28][10] = 5'd0;
    frame1[29][10] = 5'd0;
    frame1[30][10] = 5'd0;
    frame1[31][10] = 5'd0;
    frame1[0][11] = 5'd0;
    frame1[1][11] = 5'd0;
    frame1[2][11] = 5'd0;
    frame1[3][11] = 5'd0;
    frame1[4][11] = 5'd0;
    frame1[5][11] = 5'd0;
    frame1[6][11] = 5'd0;
    frame1[7][11] = 5'd0;
    frame1[8][11] = 5'd0;
    frame1[9][11] = 5'd0;
    frame1[10][11] = 5'd0;
    frame1[11][11] = 5'd0;
    frame1[12][11] = 5'd0;
    frame1[13][11] = 5'd0;
    frame1[14][11] = 5'd0;
    frame1[15][11] = 5'd0;
    frame1[16][11] = 5'd0;
    frame1[17][11] = 5'd0;
    frame1[18][11] = 5'd0;
    frame1[19][11] = 5'd0;
    frame1[20][11] = 5'd0;
    frame1[21][11] = 5'd0;
    frame1[22][11] = 5'd0;
    frame1[23][11] = 5'd0;
    frame1[24][11] = 5'd0;
    frame1[25][11] = 5'd0;
    frame1[26][11] = 5'd0;
    frame1[27][11] = 5'd0;
    frame1[28][11] = 5'd0;
    frame1[29][11] = 5'd0;
    frame1[30][11] = 5'd0;
    frame1[31][11] = 5'd0;
    frame1[0][12] = 5'd0;
    frame1[1][12] = 5'd0;
    frame1[2][12] = 5'd0;
    frame1[3][12] = 5'd0;
    frame1[4][12] = 5'd0;
    frame1[5][12] = 5'd0;
    frame1[6][12] = 5'd0;
    frame1[7][12] = 5'd0;
    frame1[8][12] = 5'd0;
    frame1[9][12] = 5'd0;
    frame1[10][12] = 5'd0;
    frame1[11][12] = 5'd0;
    frame1[12][12] = 5'd0;
    frame1[13][12] = 5'd0;
    frame1[14][12] = 5'd0;
    frame1[15][12] = 5'd0;
    frame1[16][12] = 5'd0;
    frame1[17][12] = 5'd0;
    frame1[18][12] = 5'd0;
    frame1[19][12] = 5'd0;
    frame1[20][12] = 5'd0;
    frame1[21][12] = 5'd0;
    frame1[22][12] = 5'd0;
    frame1[23][12] = 5'd0;
    frame1[24][12] = 5'd0;
    frame1[25][12] = 5'd0;
    frame1[26][12] = 5'd0;
    frame1[27][12] = 5'd0;
    frame1[28][12] = 5'd0;
    frame1[29][12] = 5'd0;
    frame1[30][12] = 5'd0;
    frame1[31][12] = 5'd0;
    frame1[0][13] = 5'd0;
    frame1[1][13] = 5'd0;
    frame1[2][13] = 5'd0;
    frame1[3][13] = 5'd0;
    frame1[4][13] = 5'd0;
    frame1[5][13] = 5'd0;
    frame1[6][13] = 5'd0;
    frame1[7][13] = 5'd0;
    frame1[8][13] = 5'd0;
    frame1[9][13] = 5'd0;
    frame1[10][13] = 5'd0;
    frame1[11][13] = 5'd0;
    frame1[12][13] = 5'd0;
    frame1[13][13] = 5'd0;
    frame1[14][13] = 5'd0;
    frame1[15][13] = 5'd0;
    frame1[16][13] = 5'd0;
    frame1[17][13] = 5'd0;
    frame1[18][13] = 5'd0;
    frame1[19][13] = 5'd0;
    frame1[20][13] = 5'd0;
    frame1[21][13] = 5'd0;
    frame1[22][13] = 5'd0;
    frame1[23][13] = 5'd0;
    frame1[24][13] = 5'd0;
    frame1[25][13] = 5'd0;
    frame1[26][13] = 5'd0;
    frame1[27][13] = 5'd0;
    frame1[28][13] = 5'd0;
    frame1[29][13] = 5'd0;
    frame1[30][13] = 5'd0;
    frame1[31][13] = 5'd0;
    frame1[0][14] = 5'd0;
    frame1[1][14] = 5'd0;
    frame1[2][14] = 5'd0;
    frame1[3][14] = 5'd0;
    frame1[4][14] = 5'd0;
    frame1[5][14] = 5'd0;
    frame1[6][14] = 5'd0;
    frame1[7][14] = 5'd0;
    frame1[8][14] = 5'd0;
    frame1[9][14] = 5'd0;
    frame1[10][14] = 5'd0;
    frame1[11][14] = 5'd0;
    frame1[12][14] = 5'd0;
    frame1[13][14] = 5'd0;
    frame1[14][14] = 5'd0;
    frame1[15][14] = 5'd0;
    frame1[16][14] = 5'd0;
    frame1[17][14] = 5'd0;
    frame1[18][14] = 5'd0;
    frame1[19][14] = 5'd0;
    frame1[20][14] = 5'd0;
    frame1[21][14] = 5'd0;
    frame1[22][14] = 5'd0;
    frame1[23][14] = 5'd0;
    frame1[24][14] = 5'd0;
    frame1[25][14] = 5'd0;
    frame1[26][14] = 5'd0;
    frame1[27][14] = 5'd0;
    frame1[28][14] = 5'd0;
    frame1[29][14] = 5'd0;
    frame1[30][14] = 5'd0;
    frame1[31][14] = 5'd0;
    frame1[0][15] = 5'd0;
    frame1[1][15] = 5'd0;
    frame1[2][15] = 5'd0;
    frame1[3][15] = 5'd0;
    frame1[4][15] = 5'd0;
    frame1[5][15] = 5'd0;
    frame1[6][15] = 5'd0;
    frame1[7][15] = 5'd0;
    frame1[8][15] = 5'd0;
    frame1[9][15] = 5'd0;
    frame1[10][15] = 5'd0;
    frame1[11][15] = 5'd0;
    frame1[12][15] = 5'd0;
    frame1[13][15] = 5'd0;
    frame1[14][15] = 5'd0;
    frame1[15][15] = 5'd0;
    frame1[16][15] = 5'd0;
    frame1[17][15] = 5'd0;
    frame1[18][15] = 5'd0;
    frame1[19][15] = 5'd0;
    frame1[20][15] = 5'd0;
    frame1[21][15] = 5'd0;
    frame1[22][15] = 5'd0;
    frame1[23][15] = 5'd0;
    frame1[24][15] = 5'd0;
    frame1[25][15] = 5'd0;
    frame1[26][15] = 5'd0;
    frame1[27][15] = 5'd0;
    frame1[28][15] = 5'd0;
    frame1[29][15] = 5'd0;
    frame1[30][15] = 5'd0;
    frame1[31][15] = 5'd0;
    frame1[0][16] = 5'd0;
    frame1[1][16] = 5'd0;
    frame1[2][16] = 5'd0;
    frame1[3][16] = 5'd0;
    frame1[4][16] = 5'd0;
    frame1[5][16] = 5'd0;
    frame1[6][16] = 5'd0;
    frame1[7][16] = 5'd0;
    frame1[8][16] = 5'd0;
    frame1[9][16] = 5'd0;
    frame1[10][16] = 5'd0;
    frame1[11][16] = 5'd0;
    frame1[12][16] = 5'd0;
    frame1[13][16] = 5'd0;
    frame1[14][16] = 5'd0;
    frame1[15][16] = 5'd0;
    frame1[16][16] = 5'd0;
    frame1[17][16] = 5'd0;
    frame1[18][16] = 5'd0;
    frame1[19][16] = 5'd0;
    frame1[20][16] = 5'd0;
    frame1[21][16] = 5'd0;
    frame1[22][16] = 5'd0;
    frame1[23][16] = 5'd0;
    frame1[24][16] = 5'd0;
    frame1[25][16] = 5'd0;
    frame1[26][16] = 5'd0;
    frame1[27][16] = 5'd0;
    frame1[28][16] = 5'd0;
    frame1[29][16] = 5'd0;
    frame1[30][16] = 5'd0;
    frame1[31][16] = 5'd0;
    frame1[0][17] = 5'd0;
    frame1[1][17] = 5'd0;
    frame1[2][17] = 5'd0;
    frame1[3][17] = 5'd0;
    frame1[4][17] = 5'd0;
    frame1[5][17] = 5'd0;
    frame1[6][17] = 5'd0;
    frame1[7][17] = 5'd0;
    frame1[8][17] = 5'd0;
    frame1[9][17] = 5'd0;
    frame1[10][17] = 5'd0;
    frame1[11][17] = 5'd0;
    frame1[12][17] = 5'd0;
    frame1[13][17] = 5'd0;
    frame1[14][17] = 5'd0;
    frame1[15][17] = 5'd0;
    frame1[16][17] = 5'd0;
    frame1[17][17] = 5'd0;
    frame1[18][17] = 5'd0;
    frame1[19][17] = 5'd0;
    frame1[20][17] = 5'd0;
    frame1[21][17] = 5'd0;
    frame1[22][17] = 5'd0;
    frame1[23][17] = 5'd0;
    frame1[24][17] = 5'd0;
    frame1[25][17] = 5'd0;
    frame1[26][17] = 5'd0;
    frame1[27][17] = 5'd0;
    frame1[28][17] = 5'd0;
    frame1[29][17] = 5'd0;
    frame1[30][17] = 5'd0;
    frame1[31][17] = 5'd0;
    frame1[0][18] = 5'd0;
    frame1[1][18] = 5'd0;
    frame1[2][18] = 5'd0;
    frame1[3][18] = 5'd0;
    frame1[4][18] = 5'd0;
    frame1[5][18] = 5'd0;
    frame1[6][18] = 5'd0;
    frame1[7][18] = 5'd0;
    frame1[8][18] = 5'd0;
    frame1[9][18] = 5'd0;
    frame1[10][18] = 5'd0;
    frame1[11][18] = 5'd0;
    frame1[12][18] = 5'd0;
    frame1[13][18] = 5'd0;
    frame1[14][18] = 5'd0;
    frame1[15][18] = 5'd0;
    frame1[16][18] = 5'd0;
    frame1[17][18] = 5'd0;
    frame1[18][18] = 5'd0;
    frame1[19][18] = 5'd0;
    frame1[20][18] = 5'd0;
    frame1[21][18] = 5'd0;
    frame1[22][18] = 5'd0;
    frame1[23][18] = 5'd0;
    frame1[24][18] = 5'd0;
    frame1[25][18] = 5'd0;
    frame1[26][18] = 5'd0;
    frame1[27][18] = 5'd0;
    frame1[28][18] = 5'd0;
    frame1[29][18] = 5'd0;
    frame1[30][18] = 5'd0;
    frame1[31][18] = 5'd0;
    frame1[0][19] = 5'd0;
    frame1[1][19] = 5'd0;
    frame1[2][19] = 5'd0;
    frame1[3][19] = 5'd0;
    frame1[4][19] = 5'd0;
    frame1[5][19] = 5'd0;
    frame1[6][19] = 5'd0;
    frame1[7][19] = 5'd0;
    frame1[8][19] = 5'd0;
    frame1[9][19] = 5'd0;
    frame1[10][19] = 5'd0;
    frame1[11][19] = 5'd0;
    frame1[12][19] = 5'd0;
    frame1[13][19] = 5'd0;
    frame1[14][19] = 5'd0;
    frame1[15][19] = 5'd0;
    frame1[16][19] = 5'd0;
    frame1[17][19] = 5'd0;
    frame1[18][19] = 5'd0;
    frame1[19][19] = 5'd0;
    frame1[20][19] = 5'd0;
    frame1[21][19] = 5'd0;
    frame1[22][19] = 5'd0;
    frame1[23][19] = 5'd0;
    frame1[24][19] = 5'd0;
    frame1[25][19] = 5'd0;
    frame1[26][19] = 5'd0;
    frame1[27][19] = 5'd0;
    frame1[28][19] = 5'd0;
    frame1[29][19] = 5'd0;
    frame1[30][19] = 5'd0;
    frame1[31][19] = 5'd0;
    frame1[0][20] = 5'd0;
    frame1[1][20] = 5'd0;
    frame1[2][20] = 5'd0;
    frame1[3][20] = 5'd0;
    frame1[4][20] = 5'd0;
    frame1[5][20] = 5'd0;
    frame1[6][20] = 5'd0;
    frame1[7][20] = 5'd0;
    frame1[8][20] = 5'd0;
    frame1[9][20] = 5'd0;
    frame1[10][20] = 5'd0;
    frame1[11][20] = 5'd0;
    frame1[12][20] = 5'd0;
    frame1[13][20] = 5'd0;
    frame1[14][20] = 5'd0;
    frame1[15][20] = 5'd0;
    frame1[16][20] = 5'd0;
    frame1[17][20] = 5'd0;
    frame1[18][20] = 5'd0;
    frame1[19][20] = 5'd0;
    frame1[20][20] = 5'd0;
    frame1[21][20] = 5'd0;
    frame1[22][20] = 5'd0;
    frame1[23][20] = 5'd0;
    frame1[24][20] = 5'd0;
    frame1[25][20] = 5'd0;
    frame1[26][20] = 5'd0;
    frame1[27][20] = 5'd0;
    frame1[28][20] = 5'd0;
    frame1[29][20] = 5'd0;
    frame1[30][20] = 5'd0;
    frame1[31][20] = 5'd0;
    frame1[0][21] = 5'd0;
    frame1[1][21] = 5'd0;
    frame1[2][21] = 5'd0;
    frame1[3][21] = 5'd0;
    frame1[4][21] = 5'd0;
    frame1[5][21] = 5'd0;
    frame1[6][21] = 5'd0;
    frame1[7][21] = 5'd0;
    frame1[8][21] = 5'd0;
    frame1[9][21] = 5'd0;
    frame1[10][21] = 5'd0;
    frame1[11][21] = 5'd0;
    frame1[12][21] = 5'd0;
    frame1[13][21] = 5'd0;
    frame1[14][21] = 5'd0;
    frame1[15][21] = 5'd0;
    frame1[16][21] = 5'd0;
    frame1[17][21] = 5'd0;
    frame1[18][21] = 5'd0;
    frame1[19][21] = 5'd0;
    frame1[20][21] = 5'd0;
    frame1[21][21] = 5'd0;
    frame1[22][21] = 5'd0;
    frame1[23][21] = 5'd0;
    frame1[24][21] = 5'd0;
    frame1[25][21] = 5'd0;
    frame1[26][21] = 5'd0;
    frame1[27][21] = 5'd0;
    frame1[28][21] = 5'd0;
    frame1[29][21] = 5'd0;
    frame1[30][21] = 5'd0;
    frame1[31][21] = 5'd0;
    frame1[0][22] = 5'd0;
    frame1[1][22] = 5'd0;
    frame1[2][22] = 5'd0;
    frame1[3][22] = 5'd0;
    frame1[4][22] = 5'd0;
    frame1[5][22] = 5'd0;
    frame1[6][22] = 5'd0;
    frame1[7][22] = 5'd0;
    frame1[8][22] = 5'd0;
    frame1[9][22] = 5'd0;
    frame1[10][22] = 5'd0;
    frame1[11][22] = 5'd0;
    frame1[12][22] = 5'd0;
    frame1[13][22] = 5'd0;
    frame1[14][22] = 5'd0;
    frame1[15][22] = 5'd0;
    frame1[16][22] = 5'd0;
    frame1[17][22] = 5'd0;
    frame1[18][22] = 5'd0;
    frame1[19][22] = 5'd0;
    frame1[20][22] = 5'd0;
    frame1[21][22] = 5'd0;
    frame1[22][22] = 5'd0;
    frame1[23][22] = 5'd0;
    frame1[24][22] = 5'd0;
    frame1[25][22] = 5'd0;
    frame1[26][22] = 5'd0;
    frame1[27][22] = 5'd0;
    frame1[28][22] = 5'd0;
    frame1[29][22] = 5'd0;
    frame1[30][22] = 5'd0;
    frame1[31][22] = 5'd0;
    frame1[0][23] = 5'd0;
    frame1[1][23] = 5'd0;
    frame1[2][23] = 5'd0;
    frame1[3][23] = 5'd0;
    frame1[4][23] = 5'd0;
    frame1[5][23] = 5'd0;
    frame1[6][23] = 5'd0;
    frame1[7][23] = 5'd0;
    frame1[8][23] = 5'd0;
    frame1[9][23] = 5'd0;
    frame1[10][23] = 5'd0;
    frame1[11][23] = 5'd0;
    frame1[12][23] = 5'd0;
    frame1[13][23] = 5'd0;
    frame1[14][23] = 5'd0;
    frame1[15][23] = 5'd0;
    frame1[16][23] = 5'd0;
    frame1[17][23] = 5'd0;
    frame1[18][23] = 5'd0;
    frame1[19][23] = 5'd0;
    frame1[20][23] = 5'd0;
    frame1[21][23] = 5'd0;
    frame1[22][23] = 5'd0;
    frame1[23][23] = 5'd0;
    frame1[24][23] = 5'd0;
    frame1[25][23] = 5'd0;
    frame1[26][23] = 5'd0;
    frame1[27][23] = 5'd0;
    frame1[28][23] = 5'd0;
    frame1[29][23] = 5'd0;
    frame1[30][23] = 5'd0;
    frame1[31][23] = 5'd0;
    frame1[0][24] = 5'd0;
    frame1[1][24] = 5'd0;
    frame1[2][24] = 5'd0;
    frame1[3][24] = 5'd0;
    frame1[4][24] = 5'd0;
    frame1[5][24] = 5'd0;
    frame1[6][24] = 5'd0;
    frame1[7][24] = 5'd0;
    frame1[8][24] = 5'd0;
    frame1[9][24] = 5'd0;
    frame1[10][24] = 5'd0;
    frame1[11][24] = 5'd0;
    frame1[12][24] = 5'd0;
    frame1[13][24] = 5'd0;
    frame1[14][24] = 5'd0;
    frame1[15][24] = 5'd0;
    frame1[16][24] = 5'd15;
    frame1[17][24] = 5'd3;
    frame1[18][24] = 5'd3;
    frame1[19][24] = 5'd3;
    frame1[20][24] = 5'd3;
    frame1[21][24] = 5'd3;
    frame1[22][24] = 5'd3;
    frame1[23][24] = 5'd3;
    frame1[24][24] = 5'd3;
    frame1[25][24] = 5'd0;
    frame1[26][24] = 5'd0;
    frame1[27][24] = 5'd0;
    frame1[28][24] = 5'd0;
    frame1[29][24] = 5'd0;
    frame1[30][24] = 5'd0;
    frame1[31][24] = 5'd0;
    frame1[0][25] = 5'd0;
    frame1[1][25] = 5'd0;
    frame1[2][25] = 5'd0;
    frame1[3][25] = 5'd0;
    frame1[4][25] = 5'd0;
    frame1[5][25] = 5'd0;
    frame1[6][25] = 5'd0;
    frame1[7][25] = 5'd0;
    frame1[8][25] = 5'd0;
    frame1[9][25] = 5'd0;
    frame1[10][25] = 5'd0;
    frame1[11][25] = 5'd0;
    frame1[12][25] = 5'd0;
    frame1[13][25] = 5'd0;
    frame1[14][25] = 5'd0;
    frame1[15][25] = 5'd0;
    frame1[16][25] = 5'd22;
    frame1[17][25] = 5'd9;
    frame1[18][25] = 5'd9;
    frame1[19][25] = 5'd9;
    frame1[20][25] = 5'd9;
    frame1[21][25] = 5'd9;
    frame1[22][25] = 5'd9;
    frame1[23][25] = 5'd9;
    frame1[24][25] = 5'd9;
    frame1[25][25] = 5'd14;
    frame1[26][25] = 5'd0;
    frame1[27][25] = 5'd0;
    frame1[28][25] = 5'd0;
    frame1[29][25] = 5'd0;
    frame1[30][25] = 5'd0;
    frame1[31][25] = 5'd0;
    frame1[0][26] = 5'd0;
    frame1[1][26] = 5'd0;
    frame1[2][26] = 5'd0;
    frame1[3][26] = 5'd0;
    frame1[4][26] = 5'd0;
    frame1[5][26] = 5'd0;
    frame1[6][26] = 5'd0;
    frame1[7][26] = 5'd0;
    frame1[8][26] = 5'd0;
    frame1[9][26] = 5'd0;
    frame1[10][26] = 5'd0;
    frame1[11][26] = 5'd0;
    frame1[12][26] = 5'd0;
    frame1[13][26] = 5'd0;
    frame1[14][26] = 5'd0;
    frame1[15][26] = 5'd15;
    frame1[16][26] = 5'd9;
    frame1[17][26] = 5'd13;
    frame1[18][26] = 5'd1;
    frame1[19][26] = 5'd1;
    frame1[20][26] = 5'd1;
    frame1[21][26] = 5'd1;
    frame1[22][26] = 5'd1;
    frame1[23][26] = 5'd1;
    frame1[24][26] = 5'd9;
    frame1[25][26] = 5'd16;
    frame1[26][26] = 5'd0;
    frame1[27][26] = 5'd0;
    frame1[28][26] = 5'd0;
    frame1[29][26] = 5'd0;
    frame1[30][26] = 5'd0;
    frame1[31][26] = 5'd0;
    frame1[0][27] = 5'd0;
    frame1[1][27] = 5'd0;
    frame1[2][27] = 5'd0;
    frame1[3][27] = 5'd0;
    frame1[4][27] = 5'd5;
    frame1[5][27] = 5'd5;
    frame1[6][27] = 5'd5;
    frame1[7][27] = 5'd5;
    frame1[8][27] = 5'd0;
    frame1[9][27] = 5'd0;
    frame1[10][27] = 5'd0;
    frame1[11][27] = 5'd0;
    frame1[12][27] = 5'd5;
    frame1[13][27] = 5'd5;
    frame1[14][27] = 5'd5;
    frame1[15][27] = 5'd21;
    frame1[16][27] = 5'd9;
    frame1[17][27] = 5'd1;
    frame1[18][27] = 5'd1;
    frame1[19][27] = 5'd1;
    frame1[20][27] = 5'd17;
    frame1[21][27] = 5'd19;
    frame1[22][27] = 5'd1;
    frame1[23][27] = 5'd1;
    frame1[24][27] = 5'd31;
    frame1[25][27] = 5'd16;
    frame1[26][27] = 5'd0;
    frame1[27][27] = 5'd0;
    frame1[28][27] = 5'd0;
    frame1[29][27] = 5'd0;
    frame1[30][27] = 5'd0;
    frame1[31][27] = 5'd0;
    frame1[0][28] = 5'd0;
    frame1[1][28] = 5'd0;
    frame1[2][28] = 5'd0;
    frame1[3][28] = 5'd0;
    frame1[4][28] = 5'd5;
    frame1[5][28] = 5'd5;
    frame1[6][28] = 5'd5;
    frame1[7][28] = 5'd5;
    frame1[8][28] = 5'd0;
    frame1[9][28] = 5'd0;
    frame1[10][28] = 5'd0;
    frame1[11][28] = 5'd0;
    frame1[12][28] = 5'd5;
    frame1[13][28] = 5'd5;
    frame1[14][28] = 5'd5;
    frame1[15][28] = 5'd21;
    frame1[16][28] = 5'd13;
    frame1[17][28] = 5'd19;
    frame1[18][28] = 5'd1;
    frame1[19][28] = 5'd1;
    frame1[20][28] = 5'd1;
    frame1[21][28] = 5'd1;
    frame1[22][28] = 5'd1;
    frame1[23][28] = 5'd1;
    frame1[24][28] = 5'd1;
    frame1[25][28] = 5'd16;
    frame1[26][28] = 5'd0;
    frame1[27][28] = 5'd0;
    frame1[28][28] = 5'd0;
    frame1[29][28] = 5'd0;
    frame1[30][28] = 5'd0;
    frame1[31][28] = 5'd0;
    frame1[0][29] = 5'd0;
    frame1[1][29] = 5'd0;
    frame1[2][29] = 5'd0;
    frame1[3][29] = 5'd0;
    frame1[4][29] = 5'd4;
    frame1[5][29] = 5'd4;
    frame1[6][29] = 5'd4;
    frame1[7][29] = 5'd4;
    frame1[8][29] = 5'd5;
    frame1[9][29] = 5'd5;
    frame1[10][29] = 5'd5;
    frame1[11][29] = 5'd5;
    frame1[12][29] = 5'd4;
    frame1[13][29] = 5'd4;
    frame1[14][29] = 5'd4;
    frame1[15][29] = 5'd28;
    frame1[16][29] = 5'd13;
    frame1[17][29] = 5'd1;
    frame1[18][29] = 5'd1;
    frame1[19][29] = 5'd1;
    frame1[20][29] = 5'd1;
    frame1[21][29] = 5'd1;
    frame1[22][29] = 5'd3;
    frame1[23][29] = 5'd19;
    frame1[24][29] = 5'd1;
    frame1[25][29] = 5'd16;
    frame1[26][29] = 5'd0;
    frame1[27][29] = 5'd3;
    frame1[28][29] = 5'd0;
    frame1[29][29] = 5'd0;
    frame1[30][29] = 5'd0;
    frame1[31][29] = 5'd0;
    frame1[0][30] = 5'd0;
    frame1[1][30] = 5'd0;
    frame1[2][30] = 5'd0;
    frame1[3][30] = 5'd0;
    frame1[4][30] = 5'd4;
    frame1[5][30] = 5'd4;
    frame1[6][30] = 5'd4;
    frame1[7][30] = 5'd4;
    frame1[8][30] = 5'd5;
    frame1[9][30] = 5'd5;
    frame1[10][30] = 5'd5;
    frame1[11][30] = 5'd5;
    frame1[12][30] = 5'd4;
    frame1[13][30] = 5'd4;
    frame1[14][30] = 5'd4;
    frame1[15][30] = 5'd28;
    frame1[16][30] = 5'd13;
    frame1[17][30] = 5'd1;
    frame1[18][30] = 5'd1;
    frame1[19][30] = 5'd1;
    frame1[20][30] = 5'd1;
    frame1[21][30] = 5'd18;
    frame1[22][30] = 5'd11;
    frame1[23][30] = 5'd1;
    frame1[24][30] = 5'd1;
    frame1[25][30] = 5'd16;
    frame1[26][30] = 5'd15;
    frame1[27][30] = 5'd2;
    frame1[28][30] = 5'd14;
    frame1[29][30] = 5'd0;
    frame1[30][30] = 5'd0;
    frame1[31][30] = 5'd0;
    frame1[0][31] = 5'd0;
    frame1[1][31] = 5'd0;
    frame1[2][31] = 5'd0;
    frame1[3][31] = 5'd0;
    frame1[4][31] = 5'd6;
    frame1[5][31] = 5'd6;
    frame1[6][31] = 5'd6;
    frame1[7][31] = 5'd6;
    frame1[8][31] = 5'd4;
    frame1[9][31] = 5'd4;
    frame1[10][31] = 5'd4;
    frame1[11][31] = 5'd4;
    frame1[12][31] = 5'd6;
    frame1[13][31] = 5'd6;
    frame1[14][31] = 5'd6;
    frame1[15][31] = 5'd23;
    frame1[16][31] = 5'd13;
    frame1[17][31] = 5'd1;
    frame1[18][31] = 5'd1;
    frame1[19][31] = 5'd19;
    frame1[20][31] = 5'd1;
    frame1[21][31] = 5'd18;
    frame1[22][31] = 5'd2;
    frame1[23][31] = 5'd3;
    frame1[24][31] = 5'd1;
    frame1[25][31] = 5'd16;
    frame1[26][31] = 5'd12;
    frame1[27][31] = 5'd2;
    frame1[28][31] = 5'd14;
    frame1[29][31] = 5'd0;
    frame1[30][31] = 5'd0;
    frame1[31][31] = 5'd0;
    frame1[0][32] = 5'd0;
    frame1[1][32] = 5'd0;
    frame1[2][32] = 5'd0;
    frame1[3][32] = 5'd0;
    frame1[4][32] = 5'd6;
    frame1[5][32] = 5'd6;
    frame1[6][32] = 5'd6;
    frame1[7][32] = 5'd6;
    frame1[8][32] = 5'd4;
    frame1[9][32] = 5'd4;
    frame1[10][32] = 5'd4;
    frame1[11][32] = 5'd4;
    frame1[12][32] = 5'd6;
    frame1[13][32] = 5'd6;
    frame1[14][32] = 5'd6;
    frame1[15][32] = 5'd23;
    frame1[16][32] = 5'd13;
    frame1[17][32] = 5'd1;
    frame1[18][32] = 5'd1;
    frame1[19][32] = 5'd1;
    frame1[20][32] = 5'd1;
    frame1[21][32] = 5'd18;
    frame1[22][32] = 5'd2;
    frame1[23][32] = 5'd2;
    frame1[24][32] = 5'd3;
    frame1[25][32] = 5'd3;
    frame1[26][32] = 5'd2;
    frame1[27][32] = 5'd2;
    frame1[28][32] = 5'd14;
    frame1[29][32] = 5'd0;
    frame1[30][32] = 5'd0;
    frame1[31][32] = 5'd0;
    frame1[0][33] = 5'd0;
    frame1[1][33] = 5'd0;
    frame1[2][33] = 5'd0;
    frame1[3][33] = 5'd0;
    frame1[4][33] = 5'd7;
    frame1[5][33] = 5'd7;
    frame1[6][33] = 5'd7;
    frame1[7][33] = 5'd7;
    frame1[8][33] = 5'd6;
    frame1[9][33] = 5'd6;
    frame1[10][33] = 5'd6;
    frame1[11][33] = 5'd6;
    frame1[12][33] = 5'd7;
    frame1[13][33] = 5'd7;
    frame1[14][33] = 5'd7;
    frame1[15][33] = 5'd24;
    frame1[16][33] = 5'd13;
    frame1[17][33] = 5'd1;
    frame1[18][33] = 5'd17;
    frame1[19][33] = 5'd1;
    frame1[20][33] = 5'd1;
    frame1[21][33] = 5'd18;
    frame1[22][33] = 5'd2;
    frame1[23][33] = 5'd2;
    frame1[24][33] = 5'd2;
    frame1[25][33] = 5'd2;
    frame1[26][33] = 5'd2;
    frame1[27][33] = 5'd2;
    frame1[28][33] = 5'd14;
    frame1[29][33] = 5'd0;
    frame1[30][33] = 5'd0;
    frame1[31][33] = 5'd0;
    frame1[0][34] = 5'd0;
    frame1[1][34] = 5'd0;
    frame1[2][34] = 5'd0;
    frame1[3][34] = 5'd0;
    frame1[4][34] = 5'd7;
    frame1[5][34] = 5'd7;
    frame1[6][34] = 5'd7;
    frame1[7][34] = 5'd7;
    frame1[8][34] = 5'd6;
    frame1[9][34] = 5'd6;
    frame1[10][34] = 5'd6;
    frame1[11][34] = 5'd6;
    frame1[12][34] = 5'd7;
    frame1[13][34] = 5'd7;
    frame1[14][34] = 5'd7;
    frame1[15][34] = 5'd3;
    frame1[16][34] = 5'd13;
    frame1[17][34] = 5'd1;
    frame1[18][34] = 5'd1;
    frame1[19][34] = 5'd1;
    frame1[20][34] = 5'd17;
    frame1[21][34] = 5'd12;
    frame1[22][34] = 5'd2;
    frame1[23][34] = 5'd2;
    frame1[24][34] = 5'd2;
    frame1[25][34] = 5'd2;
    frame1[26][34] = 5'd2;
    frame1[27][34] = 5'd2;
    frame1[28][34] = 5'd11;
    frame1[29][34] = 5'd0;
    frame1[30][34] = 5'd0;
    frame1[31][34] = 5'd0;
    frame1[0][35] = 5'd0;
    frame1[1][35] = 5'd0;
    frame1[2][35] = 5'd0;
    frame1[3][35] = 5'd0;
    frame1[4][35] = 5'd10;
    frame1[5][35] = 5'd10;
    frame1[6][35] = 5'd10;
    frame1[7][35] = 5'd10;
    frame1[8][35] = 5'd7;
    frame1[9][35] = 5'd7;
    frame1[10][35] = 5'd7;
    frame1[11][35] = 5'd7;
    frame1[12][35] = 5'd10;
    frame1[13][35] = 5'd30;
    frame1[14][35] = 5'd3;
    frame1[15][35] = 5'd3;
    frame1[16][35] = 5'd13;
    frame1[17][35] = 5'd17;
    frame1[18][35] = 5'd1;
    frame1[19][35] = 5'd1;
    frame1[20][35] = 5'd1;
    frame1[21][35] = 5'd12;
    frame1[22][35] = 5'd2;
    frame1[23][35] = 5'd20;
    frame1[24][35] = 5'd2;
    frame1[25][35] = 5'd2;
    frame1[26][35] = 5'd20;
    frame1[27][35] = 5'd2;
    frame1[28][35] = 5'd11;
    frame1[29][35] = 5'd0;
    frame1[30][35] = 5'd0;
    frame1[31][35] = 5'd0;
    frame1[0][36] = 5'd0;
    frame1[1][36] = 5'd0;
    frame1[2][36] = 5'd0;
    frame1[3][36] = 5'd0;
    frame1[4][36] = 5'd10;
    frame1[5][36] = 5'd10;
    frame1[6][36] = 5'd10;
    frame1[7][36] = 5'd10;
    frame1[8][36] = 5'd7;
    frame1[9][36] = 5'd7;
    frame1[10][36] = 5'd7;
    frame1[11][36] = 5'd7;
    frame1[12][36] = 5'd30;
    frame1[13][36] = 5'd12;
    frame1[14][36] = 5'd2;
    frame1[15][36] = 5'd11;
    frame1[16][36] = 5'd13;
    frame1[17][36] = 5'd1;
    frame1[18][36] = 5'd1;
    frame1[19][36] = 5'd1;
    frame1[20][36] = 5'd1;
    frame1[21][36] = 5'd12;
    frame1[22][36] = 5'd2;
    frame1[23][36] = 5'd3;
    frame1[24][36] = 5'd2;
    frame1[25][36] = 5'd12;
    frame1[26][36] = 5'd3;
    frame1[27][36] = 5'd2;
    frame1[28][36] = 5'd11;
    frame1[29][36] = 5'd0;
    frame1[30][36] = 5'd0;
    frame1[31][36] = 5'd0;
    frame1[0][37] = 5'd0;
    frame1[1][37] = 5'd0;
    frame1[2][37] = 5'd0;
    frame1[3][37] = 5'd0;
    frame1[4][37] = 5'd8;
    frame1[5][37] = 5'd8;
    frame1[6][37] = 5'd8;
    frame1[7][37] = 5'd8;
    frame1[8][37] = 5'd10;
    frame1[9][37] = 5'd10;
    frame1[10][37] = 5'd10;
    frame1[11][37] = 5'd10;
    frame1[12][37] = 5'd29;
    frame1[13][37] = 5'd2;
    frame1[14][37] = 5'd11;
    frame1[15][37] = 5'd3;
    frame1[16][37] = 5'd13;
    frame1[17][37] = 5'd1;
    frame1[18][37] = 5'd1;
    frame1[19][37] = 5'd17;
    frame1[20][37] = 5'd1;
    frame1[21][37] = 5'd12;
    frame1[22][37] = 5'd25;
    frame1[23][37] = 5'd2;
    frame1[24][37] = 5'd2;
    frame1[25][37] = 5'd2;
    frame1[26][37] = 5'd2;
    frame1[27][37] = 5'd27;
    frame1[28][37] = 5'd26;
    frame1[29][37] = 5'd0;
    frame1[30][37] = 5'd0;
    frame1[31][37] = 5'd0;
    frame1[0][38] = 5'd0;
    frame1[1][38] = 5'd0;
    frame1[2][38] = 5'd0;
    frame1[3][38] = 5'd0;
    frame1[4][38] = 5'd8;
    frame1[5][38] = 5'd8;
    frame1[6][38] = 5'd8;
    frame1[7][38] = 5'd8;
    frame1[8][38] = 5'd10;
    frame1[9][38] = 5'd10;
    frame1[10][38] = 5'd10;
    frame1[11][38] = 5'd10;
    frame1[12][38] = 5'd8;
    frame1[13][38] = 5'd3;
    frame1[14][38] = 5'd3;
    frame1[15][38] = 5'd29;
    frame1[16][38] = 5'd9;
    frame1[17][38] = 5'd19;
    frame1[18][38] = 5'd1;
    frame1[19][38] = 5'd1;
    frame1[20][38] = 5'd1;
    frame1[21][38] = 5'd12;
    frame1[22][38] = 5'd25;
    frame1[23][38] = 5'd11;
    frame1[24][38] = 5'd2;
    frame1[25][38] = 5'd12;
    frame1[26][38] = 5'd11;
    frame1[27][38] = 5'd27;
    frame1[28][38] = 5'd26;
    frame1[29][38] = 5'd0;
    frame1[30][38] = 5'd0;
    frame1[31][38] = 5'd0;
    frame1[0][39] = 5'd0;
    frame1[1][39] = 5'd0;
    frame1[2][39] = 5'd0;
    frame1[3][39] = 5'd0;
    frame1[4][39] = 5'd0;
    frame1[5][39] = 5'd0;
    frame1[6][39] = 5'd0;
    frame1[7][39] = 5'd0;
    frame1[8][39] = 5'd8;
    frame1[9][39] = 5'd8;
    frame1[10][39] = 5'd8;
    frame1[11][39] = 5'd8;
    frame1[12][39] = 5'd0;
    frame1[13][39] = 5'd0;
    frame1[14][39] = 5'd0;
    frame1[15][39] = 5'd15;
    frame1[16][39] = 5'd9;
    frame1[17][39] = 5'd13;
    frame1[18][39] = 5'd1;
    frame1[19][39] = 5'd1;
    frame1[20][39] = 5'd1;
    frame1[21][39] = 5'd18;
    frame1[22][39] = 5'd2;
    frame1[23][39] = 5'd11;
    frame1[24][39] = 5'd3;
    frame1[25][39] = 5'd3;
    frame1[26][39] = 5'd3;
    frame1[27][39] = 5'd2;
    frame1[28][39] = 5'd14;
    frame1[29][39] = 5'd0;
    frame1[30][39] = 5'd0;
    frame1[31][39] = 5'd0;
    frame1[0][40] = 5'd0;
    frame1[1][40] = 5'd0;
    frame1[2][40] = 5'd0;
    frame1[3][40] = 5'd0;
    frame1[4][40] = 5'd0;
    frame1[5][40] = 5'd0;
    frame1[6][40] = 5'd0;
    frame1[7][40] = 5'd0;
    frame1[8][40] = 5'd8;
    frame1[9][40] = 5'd8;
    frame1[10][40] = 5'd8;
    frame1[11][40] = 5'd8;
    frame1[12][40] = 5'd0;
    frame1[13][40] = 5'd0;
    frame1[14][40] = 5'd0;
    frame1[15][40] = 5'd15;
    frame1[16][40] = 5'd22;
    frame1[17][40] = 5'd9;
    frame1[18][40] = 5'd9;
    frame1[19][40] = 5'd9;
    frame1[20][40] = 5'd9;
    frame1[21][40] = 5'd9;
    frame1[22][40] = 5'd12;
    frame1[23][40] = 5'd2;
    frame1[24][40] = 5'd2;
    frame1[25][40] = 5'd2;
    frame1[26][40] = 5'd2;
    frame1[27][40] = 5'd11;
    frame1[28][40] = 5'd0;
    frame1[29][40] = 5'd0;
    frame1[30][40] = 5'd0;
    frame1[31][40] = 5'd0;
    frame1[0][41] = 5'd0;
    frame1[1][41] = 5'd0;
    frame1[2][41] = 5'd0;
    frame1[3][41] = 5'd0;
    frame1[4][41] = 5'd0;
    frame1[5][41] = 5'd0;
    frame1[6][41] = 5'd0;
    frame1[7][41] = 5'd0;
    frame1[8][41] = 5'd0;
    frame1[9][41] = 5'd0;
    frame1[10][41] = 5'd0;
    frame1[11][41] = 5'd0;
    frame1[12][41] = 5'd0;
    frame1[13][41] = 5'd0;
    frame1[14][41] = 5'd0;
    frame1[15][41] = 5'd12;
    frame1[16][41] = 5'd11;
    frame1[17][41] = 5'd3;
    frame1[18][41] = 5'd3;
    frame1[19][41] = 5'd3;
    frame1[20][41] = 5'd3;
    frame1[21][41] = 5'd3;
    frame1[22][41] = 5'd3;
    frame1[23][41] = 5'd3;
    frame1[24][41] = 5'd3;
    frame1[25][41] = 5'd3;
    frame1[26][41] = 5'd3;
    frame1[27][41] = 5'd14;
    frame1[28][41] = 5'd0;
    frame1[29][41] = 5'd0;
    frame1[30][41] = 5'd0;
    frame1[31][41] = 5'd0;
    frame1[0][42] = 5'd0;
    frame1[1][42] = 5'd0;
    frame1[2][42] = 5'd0;
    frame1[3][42] = 5'd0;
    frame1[4][42] = 5'd0;
    frame1[5][42] = 5'd0;
    frame1[6][42] = 5'd0;
    frame1[7][42] = 5'd0;
    frame1[8][42] = 5'd0;
    frame1[9][42] = 5'd0;
    frame1[10][42] = 5'd0;
    frame1[11][42] = 5'd0;
    frame1[12][42] = 5'd0;
    frame1[13][42] = 5'd0;
    frame1[14][42] = 5'd0;
    frame1[15][42] = 5'd12;
    frame1[16][42] = 5'd11;
    frame1[17][42] = 5'd15;
    frame1[18][42] = 5'd2;
    frame1[19][42] = 5'd14;
    frame1[20][42] = 5'd0;
    frame1[21][42] = 5'd0;
    frame1[22][42] = 5'd15;
    frame1[23][42] = 5'd2;
    frame1[24][42] = 5'd14;
    frame1[25][42] = 5'd12;
    frame1[26][42] = 5'd11;
    frame1[27][42] = 5'd0;
    frame1[28][42] = 5'd0;
    frame1[29][42] = 5'd0;
    frame1[30][42] = 5'd0;
    frame1[31][42] = 5'd0;
    frame1[0][43] = 5'd0;
    frame1[1][43] = 5'd0;
    frame1[2][43] = 5'd0;
    frame1[3][43] = 5'd0;
    frame1[4][43] = 5'd0;
    frame1[5][43] = 5'd0;
    frame1[6][43] = 5'd0;
    frame1[7][43] = 5'd0;
    frame1[8][43] = 5'd0;
    frame1[9][43] = 5'd0;
    frame1[10][43] = 5'd0;
    frame1[11][43] = 5'd0;
    frame1[12][43] = 5'd0;
    frame1[13][43] = 5'd0;
    frame1[14][43] = 5'd0;
    frame1[15][43] = 5'd3;
    frame1[16][43] = 5'd14;
    frame1[17][43] = 5'd0;
    frame1[18][43] = 5'd3;
    frame1[19][43] = 5'd14;
    frame1[20][43] = 5'd0;
    frame1[21][43] = 5'd0;
    frame1[22][43] = 5'd0;
    frame1[23][43] = 5'd3;
    frame1[24][43] = 5'd14;
    frame1[25][43] = 5'd15;
    frame1[26][43] = 5'd3;
    frame1[27][43] = 5'd0;
    frame1[28][43] = 5'd0;
    frame1[29][43] = 5'd0;
    frame1[30][43] = 5'd0;
    frame1[31][43] = 5'd0;
    frame1[0][44] = 5'd0;
    frame1[1][44] = 5'd0;
    frame1[2][44] = 5'd0;
    frame1[3][44] = 5'd0;
    frame1[4][44] = 5'd0;
    frame1[5][44] = 5'd0;
    frame1[6][44] = 5'd0;
    frame1[7][44] = 5'd0;
    frame1[8][44] = 5'd0;
    frame1[9][44] = 5'd0;
    frame1[10][44] = 5'd0;
    frame1[11][44] = 5'd0;
    frame1[12][44] = 5'd0;
    frame1[13][44] = 5'd0;
    frame1[14][44] = 5'd0;
    frame1[15][44] = 5'd0;
    frame1[16][44] = 5'd0;
    frame1[17][44] = 5'd0;
    frame1[18][44] = 5'd0;
    frame1[19][44] = 5'd0;
    frame1[20][44] = 5'd0;
    frame1[21][44] = 5'd0;
    frame1[22][44] = 5'd0;
    frame1[23][44] = 5'd0;
    frame1[24][44] = 5'd0;
    frame1[25][44] = 5'd0;
    frame1[26][44] = 5'd0;
    frame1[27][44] = 5'd0;
    frame1[28][44] = 5'd0;
    frame1[29][44] = 5'd0;
    frame1[30][44] = 5'd0;
    frame1[31][44] = 5'd0;
    frame1[0][45] = 5'd0;
    frame1[1][45] = 5'd0;
    frame1[2][45] = 5'd0;
    frame1[3][45] = 5'd0;
    frame1[4][45] = 5'd0;
    frame1[5][45] = 5'd0;
    frame1[6][45] = 5'd0;
    frame1[7][45] = 5'd0;
    frame1[8][45] = 5'd0;
    frame1[9][45] = 5'd0;
    frame1[10][45] = 5'd0;
    frame1[11][45] = 5'd0;
    frame1[12][45] = 5'd0;
    frame1[13][45] = 5'd0;
    frame1[14][45] = 5'd0;
    frame1[15][45] = 5'd0;
    frame1[16][45] = 5'd0;
    frame1[17][45] = 5'd0;
    frame1[18][45] = 5'd0;
    frame1[19][45] = 5'd0;
    frame1[20][45] = 5'd0;
    frame1[21][45] = 5'd0;
    frame1[22][45] = 5'd0;
    frame1[23][45] = 5'd0;
    frame1[24][45] = 5'd0;
    frame1[25][45] = 5'd0;
    frame1[26][45] = 5'd0;
    frame1[27][45] = 5'd0;
    frame1[28][45] = 5'd0;
    frame1[29][45] = 5'd0;
    frame1[30][45] = 5'd0;
    frame1[31][45] = 5'd0;
    frame1[0][46] = 5'd0;
    frame1[1][46] = 5'd0;
    frame1[2][46] = 5'd0;
    frame1[3][46] = 5'd0;
    frame1[4][46] = 5'd0;
    frame1[5][46] = 5'd0;
    frame1[6][46] = 5'd0;
    frame1[7][46] = 5'd0;
    frame1[8][46] = 5'd0;
    frame1[9][46] = 5'd0;
    frame1[10][46] = 5'd0;
    frame1[11][46] = 5'd0;
    frame1[12][46] = 5'd0;
    frame1[13][46] = 5'd0;
    frame1[14][46] = 5'd0;
    frame1[15][46] = 5'd0;
    frame1[16][46] = 5'd0;
    frame1[17][46] = 5'd0;
    frame1[18][46] = 5'd0;
    frame1[19][46] = 5'd0;
    frame1[20][46] = 5'd0;
    frame1[21][46] = 5'd0;
    frame1[22][46] = 5'd0;
    frame1[23][46] = 5'd0;
    frame1[24][46] = 5'd0;
    frame1[25][46] = 5'd0;
    frame1[26][46] = 5'd0;
    frame1[27][46] = 5'd0;
    frame1[28][46] = 5'd0;
    frame1[29][46] = 5'd0;
    frame1[30][46] = 5'd0;
    frame1[31][46] = 5'd0;
    frame1[0][47] = 5'd0;
    frame1[1][47] = 5'd0;
    frame1[2][47] = 5'd0;
    frame1[3][47] = 5'd0;
    frame1[4][47] = 5'd0;
    frame1[5][47] = 5'd0;
    frame1[6][47] = 5'd0;
    frame1[7][47] = 5'd0;
    frame1[8][47] = 5'd0;
    frame1[9][47] = 5'd0;
    frame1[10][47] = 5'd0;
    frame1[11][47] = 5'd0;
    frame1[12][47] = 5'd0;
    frame1[13][47] = 5'd0;
    frame1[14][47] = 5'd0;
    frame1[15][47] = 5'd0;
    frame1[16][47] = 5'd0;
    frame1[17][47] = 5'd0;
    frame1[18][47] = 5'd0;
    frame1[19][47] = 5'd0;
    frame1[20][47] = 5'd0;
    frame1[21][47] = 5'd0;
    frame1[22][47] = 5'd0;
    frame1[23][47] = 5'd0;
    frame1[24][47] = 5'd0;
    frame1[25][47] = 5'd0;
    frame1[26][47] = 5'd0;
    frame1[27][47] = 5'd0;
    frame1[28][47] = 5'd0;
    frame1[29][47] = 5'd0;
    frame1[30][47] = 5'd0;
    frame1[31][47] = 5'd0;
end

reg [5:0] palette[63:0][3:0];
initial begin
    palette[0][0] = 6'b000111;
    palette[0][1] = 6'b000111;
    palette[0][2] = 6'b000111;
    palette[0][3] = 6'b000111;
    palette[1][0] = 6'b111011;
    palette[1][1] = 6'b111011;
    palette[1][2] = 6'b111011;
    palette[1][3] = 6'b111011;
    palette[2][0] = 6'b101010;
    palette[2][1] = 6'b101010;
    palette[2][2] = 6'b101010;
    palette[2][3] = 6'b101010;
    palette[3][0] = 6'b000000;
    palette[3][1] = 6'b000000;
    palette[3][2] = 6'b000000;
    palette[3][3] = 6'b000000;
    palette[4][0] = 6'b110000;
    palette[4][1] = 6'b110000;
    palette[4][2] = 6'b110000;
    palette[4][3] = 6'b110000;
    palette[5][0] = 6'b111000;
    palette[5][1] = 6'b111000;
    palette[5][2] = 6'b111000;
    palette[5][3] = 6'b111000;
    palette[6][0] = 6'b111100;
    palette[6][1] = 6'b111100;
    palette[6][2] = 6'b111100;
    palette[6][3] = 6'b111100;
    palette[7][0] = 6'b101011;
    palette[7][1] = 6'b101011;
    palette[7][2] = 6'b101011;
    palette[7][3] = 6'b101011;
    palette[8][0] = 6'b001100;
    palette[8][1] = 6'b001100;
    palette[8][2] = 6'b001100;
    palette[8][3] = 6'b001100;
    palette[9][0] = 6'b111110;
    palette[9][1] = 6'b111011;
    palette[9][2] = 6'b111011;
    palette[9][3] = 6'b111011;
    palette[10][0] = 6'b001011;
    palette[10][1] = 6'b001011;
    palette[10][2] = 6'b001011;
    palette[10][3] = 6'b001011;
    palette[11][0] = 6'b000000;
    palette[11][1] = 6'b000111;
    palette[11][2] = 6'b000111;
    palette[11][3] = 6'b000111;
    palette[12][0] = 6'b000111;
    palette[12][1] = 6'b000111;
    palette[12][2] = 6'b000111;
    palette[12][3] = 6'b000000;
    palette[13][0] = 6'b111011;
    palette[13][1] = 6'b111011;
    palette[13][2] = 6'b000000;
    palette[13][3] = 6'b101010;
    palette[14][0] = 6'b111011;
    palette[14][1] = 6'b111011;
    palette[14][2] = 6'b111011;
    palette[14][3] = 6'b000000;
    palette[15][0] = 6'b111011;
    palette[15][1] = 6'b111011;
    palette[15][2] = 6'b111110;
    palette[15][3] = 6'b000000;
    palette[16][0] = 6'b111110;
    palette[16][1] = 6'b111110;
    palette[16][2] = 6'b111110;
    palette[16][3] = 6'b111110;
    palette[17][0] = 6'b101010;
    palette[17][1] = 6'b000000;
    palette[17][2] = 6'b000111;
    palette[17][3] = 6'b000111;
    palette[18][0] = 6'b111011;
    palette[18][1] = 6'b111011;
    palette[18][2] = 6'b111011;
    palette[18][3] = 6'b110110;
    palette[19][0] = 6'b101010;
    palette[19][1] = 6'b101010;
    palette[19][2] = 6'b101010;
    palette[19][3] = 6'b000000;
    palette[20][0] = 6'b000000;
    palette[20][1] = 6'b000000;
    palette[20][2] = 6'b000111;
    palette[20][3] = 6'b000111;
    palette[21][0] = 6'b000000;
    palette[21][1] = 6'b000000;
    palette[21][2] = 6'b000000;
    palette[21][3] = 6'b000111;
    palette[22][0] = 6'b111010;
    palette[22][1] = 6'b000000;
    palette[22][2] = 6'b000111;
    palette[22][3] = 6'b000111;
    palette[23][0] = 6'b111100;
    palette[23][1] = 6'b111100;
    palette[23][2] = 6'b111100;
    palette[23][3] = 6'b000000;
    palette[24][0] = 6'b111000;
    palette[24][1] = 6'b111000;
    palette[24][2] = 6'b111000;
    palette[24][3] = 6'b000000;
    palette[25][0] = 6'b111110;
    palette[25][1] = 6'b111011;
    palette[25][2] = 6'b111011;
    palette[25][3] = 6'b110110;
    palette[26][0] = 6'b110000;
    palette[26][1] = 6'b110000;
    palette[26][2] = 6'b110000;
    palette[26][3] = 6'b000000;
    palette[27][0] = 6'b111110;
    palette[27][1] = 6'b111110;
    palette[27][2] = 6'b111011;
    palette[27][3] = 6'b111011;
    palette[28][0] = 6'b101010;
    palette[28][1] = 6'b101010;
    palette[28][2] = 6'b000000;
    palette[28][3] = 6'b101010;
    palette[29][0] = 6'b101010;
    palette[29][1] = 6'b101010;
    palette[29][2] = 6'b000000;
    palette[29][3] = 6'b000000;
    palette[30][0] = 6'b000000;
    palette[30][1] = 6'b000000;
    palette[30][2] = 6'b101010;
    palette[30][3] = 6'b101010;
    palette[31][0] = 6'b000111;
    palette[31][1] = 6'b000111;
    palette[31][2] = 6'b000000;
    palette[31][3] = 6'b000000;
    palette[32][0] = 6'b000000;
    palette[32][1] = 6'b101010;
    palette[32][2] = 6'b101010;
    palette[32][3] = 6'b101010;
    palette[33][0] = 6'b000000;
    palette[33][1] = 6'b111110;
    palette[33][2] = 6'b111110;
    palette[33][3] = 6'b111110;
    palette[34][0] = 6'b101010;
    palette[34][1] = 6'b101010;
    palette[34][2] = 6'b000000;
    palette[34][3] = 6'b000111;
    palette[35][0] = 6'b000111;
    palette[35][1] = 6'b000111;
    palette[35][2] = 6'b000000;
    palette[35][3] = 6'b101010;
    palette[36][0] = 6'b000111;
    palette[36][1] = 6'b000000;
    palette[36][2] = 6'b101010;
    palette[36][3] = 6'b101010;
    palette[37][0] = 6'b101010;
    palette[37][1] = 6'b000000;
    palette[37][2] = 6'b000000;
    palette[37][3] = 6'b000000;
    palette[38][0] = 6'b001100;
    palette[38][1] = 6'b001100;
    palette[38][2] = 6'b001100;
    palette[38][3] = 6'b000000;
    palette[39][0] = 6'b000111;
    palette[39][1] = 6'b000000;
    palette[39][2] = 6'b000000;
    palette[39][3] = 6'b000000;
    palette[40][0] = 6'b111010;
    palette[40][1] = 6'b111010;
    palette[40][2] = 6'b101010;
    palette[40][3] = 6'b101010;
    palette[41][0] = 6'b111111;
    palette[41][1] = 6'b000000;
    palette[41][2] = 6'b101010;
    palette[41][3] = 6'b101010;
    palette[42][0] = 6'b111011;
    palette[42][1] = 6'b111110;
    palette[42][2] = 6'b111110;
    palette[42][3] = 6'b000000;
    palette[43][0] = 6'b111110;
    palette[43][1] = 6'b111011;
    palette[43][2] = 6'b110110;
    palette[43][3] = 6'b111011;
    palette[44][0] = 6'b000000;
    palette[44][1] = 6'b000000;
    palette[44][2] = 6'b111011;
    palette[44][3] = 6'b111011;
    palette[45][0] = 6'b111110;
    palette[45][1] = 6'b111110;
    palette[45][2] = 6'b000000;
    palette[45][3] = 6'b000111;
    palette[46][0] = 6'b001011;
    palette[46][1] = 6'b001011;
    palette[46][2] = 6'b000000;
    palette[46][3] = 6'b101010;
    palette[47][0] = 6'b101010;
    palette[47][1] = 6'b000000;
    palette[47][2] = 6'b111011;
    palette[47][3] = 6'b111011;
    palette[48][0] = 6'b101010;
    palette[48][1] = 6'b000000;
    palette[48][2] = 6'b101010;
    palette[48][3] = 6'b111010;
    palette[49][0] = 6'b101010;
    palette[49][1] = 6'b000000;
    palette[49][2] = 6'b000111;
    palette[49][3] = 6'b000000;
    palette[50][0] = 6'b101010;
    palette[50][1] = 6'b101010;
    palette[50][2] = 6'b101010;
    palette[50][3] = 6'b111010;
    palette[51][0] = 6'b101010;
    palette[51][1] = 6'b101010;
    palette[51][2] = 6'b111111;
    palette[51][3] = 6'b000000;
    palette[52][0] = 6'b101011;
    palette[52][1] = 6'b101011;
    palette[52][2] = 6'b101011;
    palette[52][3] = 6'b000000;
    palette[53][0] = 6'b110110;
    palette[53][1] = 6'b111011;
    palette[53][2] = 6'b111011;
    palette[53][3] = 6'b111011;
    palette[54][0] = 6'b001011;
    palette[54][1] = 6'b001011;
    palette[54][2] = 6'b001011;
    palette[54][3] = 6'b000000;
    palette[55][0] = 6'b111010;
    palette[55][1] = 6'b111010;
    palette[55][2] = 6'b101010;
    palette[55][3] = 6'b000000;
    palette[56][0] = 6'b101011;
    palette[56][1] = 6'b101011;
    palette[56][2] = 6'b000000;
    palette[56][3] = 6'b101010;
    palette[57][0] = 6'b111100;
    palette[57][1] = 6'b111100;
    palette[57][2] = 6'b000000;
    palette[57][3] = 6'b000000;
    palette[58][0] = 6'b101011;
    palette[58][1] = 6'b101011;
    palette[58][2] = 6'b000000;
    palette[58][3] = 6'b000000;
    palette[59][0] = 6'b000000;
    palette[59][1] = 6'b101010;
    palette[59][2] = 6'b101010;
    palette[59][3] = 6'b000000;
    palette[60][0] = 6'b001100;
    palette[60][1] = 6'b000000;
    palette[60][2] = 6'b101010;
    palette[60][3] = 6'b101010;
    palette[61][0] = 6'b000000;
    palette[61][1] = 6'b000111;
    palette[61][2] = 6'b000000;
    palette[61][3] = 6'b101010;
    palette[62][0] = 6'b001100;
    palette[62][1] = 6'b000000;
    palette[62][2] = 6'b101010;
    palette[62][3] = 6'b000000;
    palette[63][0] = 6'b000000;
    palette[63][1] = 6'b000000;
    palette[63][2] = 6'b101011;
    palette[63][3] = 6'b000000;
end

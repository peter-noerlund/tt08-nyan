`default_nettype none

module graphics
    #(
        parameter VGA_WIDTH = 640,
        parameter VGA_HEIGHT = 480,

        parameter H_FRONT_PORCH = 16,
        parameter H_SYNC_PULSE = 96,
        parameter H_BACK_PORCH = 48,

        parameter V_FRONT_PORCH = 10,
        parameter V_SYNC_PULSE = 2,
        parameter V_BACK_PORCH = 33
    )
    (
        input wire clk,
        input wire rst_n,

        output wire [7:0] vga_pmod
    );

    localparam X_PIXEL_BITS = $clog2(VGA_WIDTH);
    localparam Y_PIXEL_BITS = $clog2(VGA_HEIGHT);

    reg hsync;
    reg vsync;
    reg [1:0] red;
    reg [1:0] green;
    reg [1:0] blue;

    reg [X_PIXEL_BITS - 1 : 0] pixel_x;
    reg [Y_PIXEL_BITS - 1 : 0] pixel_y;

    wire [15:0] random_value;

    assign vga_pmod = {hsync, blue[1], green[1], red[1], vsync, blue[0], green[0], red[0]};

    //xorshift rng(.clk(clk), .rst_n(rst_n), .enable(1), .value(random_value));

    reg [1631 : 0] bitmap [167 : 0];
    initial begin
        bitmap[0] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[1] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[2] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[3] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[4] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[5] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[6] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[7] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[8] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[9] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[10] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[11] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[12] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[13] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[14] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[15] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[16] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[17] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[18] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[19] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[20] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[21] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[22] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[23] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[24] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[25] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[26] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[27] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[28] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[29] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[30] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[31] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[32] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[33] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[34] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[35] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[36] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[37] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[38] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[39] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[40] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[41] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[42] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[43] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[44] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[45] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[46] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[47] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[48] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[49] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[50] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[51] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[52] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[53] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[54] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[55] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[56] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[57] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[58] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[59] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[60] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[61] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[62] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[63] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111010111000000000000000000000000000000000000000000000000;
        bitmap[64] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[65] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[66] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[67] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[68] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[69] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[70] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[71] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[72] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[73] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[74] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[75] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[76] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[77] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[78] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[79] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[80] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[81] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[82] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[83] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[84] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[85] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[86] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[87] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000;
        bitmap[88] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[89] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[90] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[91] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[92] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[93] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[94] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[95] = 1632'b110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[96] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[97] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[98] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[99] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[100] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[101] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[102] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[103] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[104] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[105] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[106] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[107] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[108] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[109] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[110] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[111] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[112] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[113] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[114] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[115] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[116] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[117] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[118] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[119] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100;
        bitmap[120] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[121] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[122] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[123] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[124] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[125] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[126] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[127] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[128] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[129] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[130] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[131] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[132] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[133] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[134] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[135] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[136] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[137] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[138] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[139] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[140] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[141] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[142] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[143] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111010011010011010011010011010011010011010011010011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[144] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[145] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[146] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[147] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[148] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[149] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[150] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[151] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111110111011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[152] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[153] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[154] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[155] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[156] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[157] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[158] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[159] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011011000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[160] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[161] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[162] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[163] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[164] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[165] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[166] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
        bitmap[167] = 1632'b110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100110100;
    end
    

    always @ (posedge clk) begin
        if (!rst_n) begin
            pixel_x <= {X_PIXEL_BITS{1'b0}};
            pixel_y <= {Y_PIXEL_BITS{1'b0}};
            hsync <= 1'b1;
            vsync <= 1'b1;
            red <= 2'd0;
            green <= 2'd0;
            blue <= 2'd0;
        end else begin
            if (pixel_x == VGA_WIDTH + H_FRONT_PORCH) begin
                hsync <= 1'b1;
            end
            if (pixel_x == VGA_WIDTH + H_FRONT_PORCH + H_SYNC_PULSE) begin
                hsync <= 1'b0;
            end

            if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH) begin
                vsync <= 1'b1;
            end
            if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH + V_SYNC_PULSE) begin
                vsync <= 1'b0;
            end

            if (pixel_x == VGA_WIDTH + H_BACK_PORCH + H_SYNC_PULSE + H_BACK_PORCH - 1) begin
                pixel_x <= {X_PIXEL_BITS{1'b0}};
                if (pixel_y == VGA_HEIGHT + V_FRONT_PORCH + V_SYNC_PULSE + V_BACK_PORCH - 1) begin
                    pixel_y <= {Y_PIXEL_BITS{1'b0}};
                end else begin
                    pixel_y <= pixel_y + 1;
                end
            end else begin
                pixel_x <= pixel_x + 1;
            end

            if (pixel_x < 272 && pixel_y < 168) begin
                {blue, green, red} <= bitmap[168 - pixel_y[7:0]][(272 - pixel_x) * 6 - 1 -: 6];
            end else begin
                {red, green, blue} <= 6'b000111;
            end
            /*            
            if (pixel_x < VGA_WIDTH && pixel_y < VGA_HEIGHT) begin
                red <= random_value[1:0];
                green <= random_value[3:2];
                blue <= random_value[5:4];
            end else begin
                red <= 2'd0;
                green <= 2'd0;
                blue <= 2'd0;
            end
            */
        end
    end
endmodule
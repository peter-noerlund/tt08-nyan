reg [5:0] frame0[15:0][31:0];
initial begin
    frame0[0][0] = 6'd0;
    frame0[1][0] = 6'd0;
    frame0[2][0] = 6'd0;
    frame0[3][0] = 6'd0;
    frame0[4][0] = 6'd0;
    frame0[5][0] = 6'd0;
    frame0[6][0] = 6'd0;
    frame0[7][0] = 6'd0;
    frame0[8][0] = 6'd0;
    frame0[9][0] = 6'd0;
    frame0[10][0] = 6'd0;
    frame0[11][0] = 6'd0;
    frame0[12][0] = 6'd0;
    frame0[13][0] = 6'd0;
    frame0[14][0] = 6'd0;
    frame0[15][0] = 6'd0;
    frame0[0][1] = 6'd0;
    frame0[1][1] = 6'd0;
    frame0[2][1] = 6'd0;
    frame0[3][1] = 6'd0;
    frame0[4][1] = 6'd0;
    frame0[5][1] = 6'd0;
    frame0[6][1] = 6'd0;
    frame0[7][1] = 6'd0;
    frame0[8][1] = 6'd0;
    frame0[9][1] = 6'd0;
    frame0[10][1] = 6'd0;
    frame0[11][1] = 6'd0;
    frame0[12][1] = 6'd0;
    frame0[13][1] = 6'd0;
    frame0[14][1] = 6'd0;
    frame0[15][1] = 6'd0;
    frame0[0][2] = 6'd0;
    frame0[1][2] = 6'd0;
    frame0[2][2] = 6'd0;
    frame0[3][2] = 6'd0;
    frame0[4][2] = 6'd0;
    frame0[5][2] = 6'd0;
    frame0[6][2] = 6'd0;
    frame0[7][2] = 6'd0;
    frame0[8][2] = 6'd0;
    frame0[9][2] = 6'd0;
    frame0[10][2] = 6'd0;
    frame0[11][2] = 6'd0;
    frame0[12][2] = 6'd0;
    frame0[13][2] = 6'd0;
    frame0[14][2] = 6'd0;
    frame0[15][2] = 6'd0;
    frame0[0][3] = 6'd0;
    frame0[1][3] = 6'd0;
    frame0[2][3] = 6'd0;
    frame0[3][3] = 6'd0;
    frame0[4][3] = 6'd0;
    frame0[5][3] = 6'd0;
    frame0[6][3] = 6'd0;
    frame0[7][3] = 6'd0;
    frame0[8][3] = 6'd0;
    frame0[9][3] = 6'd0;
    frame0[10][3] = 6'd0;
    frame0[11][3] = 6'd0;
    frame0[12][3] = 6'd0;
    frame0[13][3] = 6'd0;
    frame0[14][3] = 6'd0;
    frame0[15][3] = 6'd0;
    frame0[0][4] = 6'd0;
    frame0[1][4] = 6'd0;
    frame0[2][4] = 6'd0;
    frame0[3][4] = 6'd0;
    frame0[4][4] = 6'd0;
    frame0[5][4] = 6'd0;
    frame0[6][4] = 6'd0;
    frame0[7][4] = 6'd0;
    frame0[8][4] = 6'd0;
    frame0[9][4] = 6'd0;
    frame0[10][4] = 6'd0;
    frame0[11][4] = 6'd0;
    frame0[12][4] = 6'd0;
    frame0[13][4] = 6'd0;
    frame0[14][4] = 6'd0;
    frame0[15][4] = 6'd0;
    frame0[0][5] = 6'd0;
    frame0[1][5] = 6'd0;
    frame0[2][5] = 6'd0;
    frame0[3][5] = 6'd0;
    frame0[4][5] = 6'd0;
    frame0[5][5] = 6'd0;
    frame0[6][5] = 6'd0;
    frame0[7][5] = 6'd0;
    frame0[8][5] = 6'd0;
    frame0[9][5] = 6'd0;
    frame0[10][5] = 6'd0;
    frame0[11][5] = 6'd0;
    frame0[12][5] = 6'd0;
    frame0[13][5] = 6'd0;
    frame0[14][5] = 6'd0;
    frame0[15][5] = 6'd0;
    frame0[0][6] = 6'd0;
    frame0[1][6] = 6'd0;
    frame0[2][6] = 6'd0;
    frame0[3][6] = 6'd0;
    frame0[4][6] = 6'd0;
    frame0[5][6] = 6'd0;
    frame0[6][6] = 6'd0;
    frame0[7][6] = 6'd0;
    frame0[8][6] = 6'd0;
    frame0[9][6] = 6'd0;
    frame0[10][6] = 6'd0;
    frame0[11][6] = 6'd0;
    frame0[12][6] = 6'd0;
    frame0[13][6] = 6'd0;
    frame0[14][6] = 6'd0;
    frame0[15][6] = 6'd0;
    frame0[0][7] = 6'd0;
    frame0[1][7] = 6'd0;
    frame0[2][7] = 6'd0;
    frame0[3][7] = 6'd0;
    frame0[4][7] = 6'd0;
    frame0[5][7] = 6'd0;
    frame0[6][7] = 6'd0;
    frame0[7][7] = 6'd0;
    frame0[8][7] = 6'd0;
    frame0[9][7] = 6'd0;
    frame0[10][7] = 6'd0;
    frame0[11][7] = 6'd0;
    frame0[12][7] = 6'd0;
    frame0[13][7] = 6'd0;
    frame0[14][7] = 6'd0;
    frame0[15][7] = 6'd0;
    frame0[0][8] = 6'd0;
    frame0[1][8] = 6'd0;
    frame0[2][8] = 6'd0;
    frame0[3][8] = 6'd0;
    frame0[4][8] = 6'd0;
    frame0[5][8] = 6'd0;
    frame0[6][8] = 6'd0;
    frame0[7][8] = 6'd0;
    frame0[8][8] = 6'd0;
    frame0[9][8] = 6'd0;
    frame0[10][8] = 6'd0;
    frame0[11][8] = 6'd0;
    frame0[12][8] = 6'd0;
    frame0[13][8] = 6'd0;
    frame0[14][8] = 6'd0;
    frame0[15][8] = 6'd0;
    frame0[0][9] = 6'd0;
    frame0[1][9] = 6'd0;
    frame0[2][9] = 6'd0;
    frame0[3][9] = 6'd0;
    frame0[4][9] = 6'd0;
    frame0[5][9] = 6'd0;
    frame0[6][9] = 6'd0;
    frame0[7][9] = 6'd0;
    frame0[8][9] = 6'd0;
    frame0[9][9] = 6'd0;
    frame0[10][9] = 6'd0;
    frame0[11][9] = 6'd0;
    frame0[12][9] = 6'd0;
    frame0[13][9] = 6'd0;
    frame0[14][9] = 6'd0;
    frame0[15][9] = 6'd0;
    frame0[0][10] = 6'd0;
    frame0[1][10] = 6'd0;
    frame0[2][10] = 6'd0;
    frame0[3][10] = 6'd0;
    frame0[4][10] = 6'd0;
    frame0[5][10] = 6'd0;
    frame0[6][10] = 6'd0;
    frame0[7][10] = 6'd0;
    frame0[8][10] = 6'd39;
    frame0[9][10] = 6'd3;
    frame0[10][10] = 6'd3;
    frame0[11][10] = 6'd3;
    frame0[12][10] = 6'd20;
    frame0[13][10] = 6'd0;
    frame0[14][10] = 6'd0;
    frame0[15][10] = 6'd0;
    frame0[0][11] = 6'd0;
    frame0[1][11] = 6'd0;
    frame0[2][11] = 6'd0;
    frame0[3][11] = 6'd0;
    frame0[4][11] = 6'd4;
    frame0[5][11] = 6'd4;
    frame0[6][11] = 6'd0;
    frame0[7][11] = 6'd0;
    frame0[8][11] = 6'd33;
    frame0[9][11] = 6'd16;
    frame0[10][11] = 6'd16;
    frame0[11][11] = 6'd16;
    frame0[12][11] = 6'd45;
    frame0[13][11] = 6'd0;
    frame0[14][11] = 6'd0;
    frame0[15][11] = 6'd0;
    frame0[0][12] = 6'd0;
    frame0[1][12] = 6'd0;
    frame0[2][12] = 6'd0;
    frame0[3][12] = 6'd0;
    frame0[4][12] = 6'd4;
    frame0[5][12] = 6'd4;
    frame0[6][12] = 6'd0;
    frame0[7][12] = 6'd12;
    frame0[8][12] = 6'd27;
    frame0[9][12] = 6'd1;
    frame0[10][12] = 6'd1;
    frame0[11][12] = 6'd1;
    frame0[12][12] = 6'd42;
    frame0[13][12] = 6'd0;
    frame0[14][12] = 6'd0;
    frame0[15][12] = 6'd0;
    frame0[0][13] = 6'd0;
    frame0[1][13] = 6'd0;
    frame0[2][13] = 6'd4;
    frame0[3][13] = 6'd4;
    frame0[4][13] = 6'd5;
    frame0[5][13] = 6'd5;
    frame0[6][13] = 6'd4;
    frame0[7][13] = 6'd26;
    frame0[8][13] = 6'd9;
    frame0[9][13] = 6'd1;
    frame0[10][13] = 6'd18;
    frame0[11][13] = 6'd1;
    frame0[12][13] = 6'd15;
    frame0[13][13] = 6'd0;
    frame0[14][13] = 6'd0;
    frame0[15][13] = 6'd0;
    frame0[0][14] = 6'd0;
    frame0[1][14] = 6'd0;
    frame0[2][14] = 6'd4;
    frame0[3][14] = 6'd4;
    frame0[4][14] = 6'd5;
    frame0[5][14] = 6'd5;
    frame0[6][14] = 6'd4;
    frame0[7][14] = 6'd26;
    frame0[8][14] = 6'd25;
    frame0[9][14] = 6'd1;
    frame0[10][14] = 6'd1;
    frame0[11][14] = 6'd1;
    frame0[12][14] = 6'd15;
    frame0[13][14] = 6'd0;
    frame0[14][14] = 6'd0;
    frame0[15][14] = 6'd0;
    frame0[0][15] = 6'd0;
    frame0[1][15] = 6'd0;
    frame0[2][15] = 6'd5;
    frame0[3][15] = 6'd5;
    frame0[4][15] = 6'd6;
    frame0[5][15] = 6'd6;
    frame0[6][15] = 6'd5;
    frame0[7][15] = 6'd24;
    frame0[8][15] = 6'd9;
    frame0[9][15] = 6'd1;
    frame0[10][15] = 6'd1;
    frame0[11][15] = 6'd44;
    frame0[12][15] = 6'd15;
    frame0[13][15] = 6'd31;
    frame0[14][15] = 6'd0;
    frame0[15][15] = 6'd0;
    frame0[0][16] = 6'd0;
    frame0[1][16] = 6'd0;
    frame0[2][16] = 6'd5;
    frame0[3][16] = 6'd5;
    frame0[4][16] = 6'd6;
    frame0[5][16] = 6'd6;
    frame0[6][16] = 6'd5;
    frame0[7][16] = 6'd24;
    frame0[8][16] = 6'd9;
    frame0[9][16] = 6'd1;
    frame0[10][16] = 6'd14;
    frame0[11][16] = 6'd47;
    frame0[12][16] = 6'd15;
    frame0[13][16] = 6'd36;
    frame0[14][16] = 6'd11;
    frame0[15][16] = 6'd0;
    frame0[0][17] = 6'd0;
    frame0[1][17] = 6'd0;
    frame0[2][17] = 6'd6;
    frame0[3][17] = 6'd6;
    frame0[4][17] = 6'd8;
    frame0[5][17] = 6'd8;
    frame0[6][17] = 6'd6;
    frame0[7][17] = 6'd23;
    frame0[8][17] = 6'd9;
    frame0[9][17] = 6'd18;
    frame0[10][17] = 6'd14;
    frame0[11][17] = 6'd29;
    frame0[12][17] = 6'd15;
    frame0[13][17] = 6'd32;
    frame0[14][17] = 6'd11;
    frame0[15][17] = 6'd0;
    frame0[0][18] = 6'd0;
    frame0[1][18] = 6'd0;
    frame0[2][18] = 6'd6;
    frame0[3][18] = 6'd6;
    frame0[4][18] = 6'd8;
    frame0[5][18] = 6'd8;
    frame0[6][18] = 6'd57;
    frame0[7][18] = 6'd23;
    frame0[8][18] = 6'd9;
    frame0[9][18] = 6'd1;
    frame0[10][18] = 6'd14;
    frame0[11][18] = 6'd2;
    frame0[12][18] = 6'd3;
    frame0[13][18] = 6'd2;
    frame0[14][18] = 6'd11;
    frame0[15][18] = 6'd0;
    frame0[0][19] = 6'd0;
    frame0[1][19] = 6'd0;
    frame0[2][19] = 6'd8;
    frame0[3][19] = 6'd8;
    frame0[4][19] = 6'd10;
    frame0[5][19] = 6'd10;
    frame0[6][19] = 6'd62;
    frame0[7][19] = 6'd38;
    frame0[8][19] = 6'd9;
    frame0[9][19] = 6'd53;
    frame0[10][19] = 6'd14;
    frame0[11][19] = 6'd2;
    frame0[12][19] = 6'd2;
    frame0[13][19] = 6'd2;
    frame0[14][19] = 6'd11;
    frame0[15][19] = 6'd0;
    frame0[0][20] = 6'd0;
    frame0[1][20] = 6'd0;
    frame0[2][20] = 6'd8;
    frame0[3][20] = 6'd8;
    frame0[4][20] = 6'd10;
    frame0[5][20] = 6'd10;
    frame0[6][20] = 6'd60;
    frame0[7][20] = 6'd3;
    frame0[8][20] = 6'd9;
    frame0[9][20] = 6'd1;
    frame0[10][20] = 6'd13;
    frame0[11][20] = 6'd2;
    frame0[12][20] = 6'd2;
    frame0[13][20] = 6'd2;
    frame0[14][20] = 6'd17;
    frame0[15][20] = 6'd0;
    frame0[0][21] = 6'd0;
    frame0[1][21] = 6'd0;
    frame0[2][21] = 6'd10;
    frame0[3][21] = 6'd10;
    frame0[4][21] = 6'd7;
    frame0[5][21] = 6'd7;
    frame0[6][21] = 6'd46;
    frame0[7][21] = 6'd19;
    frame0[8][21] = 6'd43;
    frame0[9][21] = 6'd1;
    frame0[10][21] = 6'd13;
    frame0[11][21] = 6'd51;
    frame0[12][21] = 6'd2;
    frame0[13][21] = 6'd41;
    frame0[14][21] = 6'd17;
    frame0[15][21] = 6'd0;
    frame0[0][22] = 6'd0;
    frame0[1][22] = 6'd0;
    frame0[2][22] = 6'd10;
    frame0[3][22] = 6'd10;
    frame0[4][22] = 6'd7;
    frame0[5][22] = 6'd7;
    frame0[6][22] = 6'd54;
    frame0[7][22] = 6'd3;
    frame0[8][22] = 6'd9;
    frame0[9][22] = 6'd18;
    frame0[10][22] = 6'd13;
    frame0[11][22] = 6'd29;
    frame0[12][22] = 6'd28;
    frame0[13][22] = 6'd30;
    frame0[14][22] = 6'd17;
    frame0[15][22] = 6'd0;
    frame0[0][23] = 6'd0;
    frame0[1][23] = 6'd0;
    frame0[2][23] = 6'd7;
    frame0[3][23] = 6'd7;
    frame0[4][23] = 6'd0;
    frame0[5][23] = 6'd0;
    frame0[6][23] = 6'd7;
    frame0[7][23] = 6'd52;
    frame0[8][23] = 6'd9;
    frame0[9][23] = 6'd1;
    frame0[10][23] = 6'd13;
    frame0[11][23] = 6'd40;
    frame0[12][23] = 6'd2;
    frame0[13][23] = 6'd50;
    frame0[14][23] = 6'd22;
    frame0[15][23] = 6'd0;
    frame0[0][24] = 6'd0;
    frame0[1][24] = 6'd0;
    frame0[2][24] = 6'd7;
    frame0[3][24] = 6'd7;
    frame0[4][24] = 6'd0;
    frame0[5][24] = 6'd0;
    frame0[6][24] = 6'd7;
    frame0[7][24] = 6'd52;
    frame0[8][24] = 6'd25;
    frame0[9][24] = 6'd1;
    frame0[10][24] = 6'd13;
    frame0[11][24] = 6'd55;
    frame0[12][24] = 6'd28;
    frame0[13][24] = 6'd48;
    frame0[14][24] = 6'd22;
    frame0[15][24] = 6'd0;
    frame0[0][25] = 6'd0;
    frame0[1][25] = 6'd0;
    frame0[2][25] = 6'd0;
    frame0[3][25] = 6'd0;
    frame0[4][25] = 6'd0;
    frame0[5][25] = 6'd0;
    frame0[6][25] = 6'd0;
    frame0[7][25] = 6'd12;
    frame0[8][25] = 6'd27;
    frame0[9][25] = 6'd1;
    frame0[10][25] = 6'd14;
    frame0[11][25] = 6'd19;
    frame0[12][25] = 6'd3;
    frame0[13][25] = 6'd30;
    frame0[14][25] = 6'd11;
    frame0[15][25] = 6'd0;
    frame0[0][26] = 6'd0;
    frame0[1][26] = 6'd0;
    frame0[2][26] = 6'd0;
    frame0[3][26] = 6'd0;
    frame0[4][26] = 6'd0;
    frame0[5][26] = 6'd0;
    frame0[6][26] = 6'd0;
    frame0[7][26] = 6'd12;
    frame0[8][26] = 6'd33;
    frame0[9][26] = 6'd16;
    frame0[10][26] = 6'd16;
    frame0[11][26] = 6'd32;
    frame0[12][26] = 6'd2;
    frame0[13][26] = 6'd19;
    frame0[14][26] = 6'd0;
    frame0[15][26] = 6'd0;
    frame0[0][27] = 6'd0;
    frame0[1][27] = 6'd0;
    frame0[2][27] = 6'd0;
    frame0[3][27] = 6'd0;
    frame0[4][27] = 6'd0;
    frame0[5][27] = 6'd0;
    frame0[6][27] = 6'd0;
    frame0[7][27] = 6'd12;
    frame0[8][27] = 6'd37;
    frame0[9][27] = 6'd3;
    frame0[10][27] = 6'd3;
    frame0[11][27] = 6'd3;
    frame0[12][27] = 6'd3;
    frame0[13][27] = 6'd21;
    frame0[14][27] = 6'd0;
    frame0[15][27] = 6'd0;
    frame0[0][28] = 6'd0;
    frame0[1][28] = 6'd0;
    frame0[2][28] = 6'd0;
    frame0[3][28] = 6'd0;
    frame0[4][28] = 6'd0;
    frame0[5][28] = 6'd0;
    frame0[6][28] = 6'd0;
    frame0[7][28] = 6'd12;
    frame0[8][28] = 6'd34;
    frame0[9][28] = 6'd59;
    frame0[10][28] = 6'd0;
    frame0[11][28] = 6'd35;
    frame0[12][28] = 6'd49;
    frame0[13][28] = 6'd34;
    frame0[14][28] = 6'd0;
    frame0[15][28] = 6'd0;
    frame0[0][29] = 6'd0;
    frame0[1][29] = 6'd0;
    frame0[2][29] = 6'd0;
    frame0[3][29] = 6'd0;
    frame0[4][29] = 6'd0;
    frame0[5][29] = 6'd0;
    frame0[6][29] = 6'd0;
    frame0[7][29] = 6'd12;
    frame0[8][29] = 6'd20;
    frame0[9][29] = 6'd39;
    frame0[10][29] = 6'd0;
    frame0[11][29] = 6'd12;
    frame0[12][29] = 6'd20;
    frame0[13][29] = 6'd21;
    frame0[14][29] = 6'd0;
    frame0[15][29] = 6'd0;
    frame0[0][30] = 6'd0;
    frame0[1][30] = 6'd0;
    frame0[2][30] = 6'd0;
    frame0[3][30] = 6'd0;
    frame0[4][30] = 6'd0;
    frame0[5][30] = 6'd0;
    frame0[6][30] = 6'd0;
    frame0[7][30] = 6'd0;
    frame0[8][30] = 6'd0;
    frame0[9][30] = 6'd0;
    frame0[10][30] = 6'd0;
    frame0[11][30] = 6'd0;
    frame0[12][30] = 6'd0;
    frame0[13][30] = 6'd0;
    frame0[14][30] = 6'd0;
    frame0[15][30] = 6'd0;
    frame0[0][31] = 6'd0;
    frame0[1][31] = 6'd0;
    frame0[2][31] = 6'd0;
    frame0[3][31] = 6'd0;
    frame0[4][31] = 6'd0;
    frame0[5][31] = 6'd0;
    frame0[6][31] = 6'd0;
    frame0[7][31] = 6'd0;
    frame0[8][31] = 6'd0;
    frame0[9][31] = 6'd0;
    frame0[10][31] = 6'd0;
    frame0[11][31] = 6'd0;
    frame0[12][31] = 6'd0;
    frame0[13][31] = 6'd0;
    frame0[14][31] = 6'd0;
    frame0[15][31] = 6'd0;
end
